XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"���-�Q(/�(3V#�
��HU��y)�x�����Q�_�\    �
$/Q�-�͓���[��
z4�D�    ���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI    �!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��R�^��E�c�i��c�X7��܄�/v��M�� �y� �Vv�ۏޕ �
�"1n����r) ��:�M�[�=}S`)9�6�%&l�G5��q����,S�c0j�d��EF��hx� )�,��+�v����f ˊ
�^�_"��藥����S��/M9�茇�:4��/@�����% �+�3��s�o��Up{��~��[���9v�5��*b��� ���*������ǆzQ�ky�c?�� �ah$!��?��m�4�>��O��Θ�G�͕��MF�zʵ��6���s,��ZP�b���W`��9G�Ϋ!�^�)҇�������&�28D:n�/4    5�R���5������ԣ�7�x�zI�.ѧ��>"�s�;�}骀s!��y&�Wl�{�����݋�0}���З�XL_�A�y"�l�Vx=�;c,6�f#��`�I�����S`�t���{�M0��?Z͸�ճ-�J��N=�ɐD�)P9��m�&��Y<(@Ț�����ÃSg��00�R3��8�\*C��y�Xv��f}��ڶt�3�h�꠹@ˆ���]�\9�#�Y�饉��y����"]z(�0���C�X'w�M�QZD���\/bn�D��/Ca&��=İa�g�_jf��e���4Q^�)�Z�E�+�Jk��j��W�z��y�IBA��r2����V�5]�J;�r���/ʱ��v 1�]���>������=�� ��l����)����g���o�r<�N+����~�Y_RXlxVHYEB     400     190�#�K|MBC�l}�A/��h�y*0�%�� ?UVA�>�Bz����k�������E�'�c���    �aė��ڰ~B��U҄r,#�����d�h�71B(���g~)+d5 �>)��dXC�k��s    �X}3������H�W�߭:t� 5\ B]�=7Vm. e�1Üv�����BIc�(ߓ��X�Bq���u�ߟiw�hNGt��o7��P�;i���b����6��cܑ�s�{C*d�J�������l ������y��;�����G��Zb05ať�D���!�?(�"�!����0�Cc��^�b+��EB��8p0z0�@�-@MV"�[��дٰ�a��:��gIl����H�Iȳ��;)�|��F�m��i_ট3�`7�XlxVHYEB     400     1c0��b{�����C�guႺ������VߪI�*~�
ER�cb��{ѭ��d��%������W~ѻ5؇�S�Nv��N&Ș&�e"[1���ނacf���~N�h�[�9�/:c`��<���2¹��Pmb�ά�ư�.v�Ѡp���o������==��ԃޭ�P��X���"��Q=��De�v{��]ݞ��w��W���HF�i��ЉRQJ��Xz��s�l3�"ڢyI8*N�.نQ0�o�*��Bo�+9o��dH\��s��|'"Ef�#�Le�>G|'\v�$r��L^e� &6�N^�����T
��w\.��d�N�vT�%��?�)��;�����V�؋y{��P5��a1К
��_C5O�P��P돈l~��J�Ŏy|B�lRͲG|;�ʥJ��A �B֥*� �?@����Mm
'�S<QłC�����66$�XlxVHYEB     400     150/�m����X�k�O\�����." nf�7���
�T@�y�L$̣^�d �*Qd���T`�*��F�B����x��r&����Go�37���͐�kp���։Q\�͵nf�����3ն���%�V`GL���.=K�sΔ�U��Q��s�k���#)� >���=T    `~aN����j�[�$�u�1Y�7�ğ�vɐ��O�����]� L�_0W?j%I�����r��x�}k˓�Z�:>�-SW��1��j�NX��� Z�Mo�漀D�����c�y��[�������4Փ@U0��,���s��*F����q�ũ��WO.)D��`���XlxVHYEB     400     170��Wx߸��z�Y��������Z�LY7�ݣr�P]╜Q�-E�|���'�#�K��Jn�Q���R~rB�e��y"� B�)��V��L"[EQ()0�Ma���|$�����}�E�����7�X[=6��#�BZ��~���}�8���fK�ɲT%�:~e�s�\����+I8��5N����&P��V�y.Q׍ߤ����������VF���.         ��s�,���dv�"Q�S5�"�8��¢|G�c]f���{�3mv��    �G�/HL��0�`ǽ��^4`��Wj��O�ͶK�VDn����$��    �=?{��6"x��aϫ����-X�e�δo���Y����hDNްj>_���j��� kik�@XlxVHYEB     400     150�)�n�H]�ע5+���Lۉ�n������R ����c�2���8jH���]�R�Öx|b�=|V�n7f!�yL��c~�L�Ͼw�l���쵦y    ��d�vP��?��<�!��q�n���4�߼�x���)*2N�F��(0�[q�9��eވ�J������̯2�D�ߙp/������wdB�;�q��i�f�9�����B�~�T�QA��{��D�Jt�MNÇ~/�`0�������K�-�B:��ğ2w��=J���u�����Ș٭��p�><�3�?�o�\B�1Ϙ�Xo�yz��A�?������'[S���Sj�W<XlxVHYEB     400     140�d��ns����PUz�wGQQG��l��`���ʐ    ��� 딄�َ g��M��*ց��eڹ;��w_Q+C����ڈp ���޸h܉���\(:|K�J1n0��"���������^�Vj�v�!�1~k7�ߓ�[&?<(�߉��.̊�D��p�g�q�1/�+����lWE^x�b<3a�5��:��%1R�W�H��fS�O�d��tP�=j��x�uh���l7�s˷g; ���s����mʛR
AX�r�9C@�Y��h���j��у_l���s�Uwۖ�³��;�3���I6)�F:}~q�<֥kXlxVHYEB     400     110y }�aq�.:/�i:������!P,��8��؍����Y�J�Wu�g2����߫#���ly�]lbB���V� ��Nu������pŹ�'���-    �����Z�Q%���8����X������lMl+�X��S�����j���'��;Y��TA"V�%Dkt8����O�ǈnyC{W��#�`K�ϙ�D.)��e�o�ȧH/�Z�m∫����[4�3b$7ƺ,"�i���U��P4/�H%W��*�����!���²XlxVHYEB     400     190|��=�����A7���fv��|�'�����)��*���Sn�Lh8��� �bR������D^��h����S�_;�@�0��F��,�e��AN?S��a�����|'$L�4ݸG7Ԯv`��M�w��yi�mL(��dK��4���Ł�
��l�R�RE�t�� �n}�DD�%������f�    �S�� .i5ó*ȣ�X��ᴲ����ܼ��zʕ�|��J�%�IE�[P@��H�s�����.�p(�%�ҹ    �z�{�Ϯ�L���-9Ъ޴U��
�����a�p6�+"���"�e�<��9�?��;���4갍ԡ����7W'��/(2���x{��J�����F��e7�L�8�t9`��U?C��AW�m���.���C=ے��%XlxVHYEB     400     160�I='��WhQtW�8,+�g1��_}pz�͏o]~�]��9���{}C�TV��AB���9�'`�x>U���ܙ����
��gb����]R ���h�����]    �L-g��\�{L=#��3�����۝�K�hg���._�B���DP�؏kc(�Rq�֤F�G5��n��B�7t�>�Uw���ȷ��"i��-�'Wa�I������g�R5Q�#�Ob�9�>��Xu"?�$��x��%%��9�55~w������g�@] ��u�7�Jw����    5�}��ix�:�#<�vS�&�J�a�}oVp��j��U9=
W��ŝD���b��z�;�c_a$HX�A1�XlxVHYEB     400     130�zto�/F����U.�̤SI�x�y7%��"Sb�;���&*>��yF�G
�`͵°��r�4������6�գu���Q�:��0d%N-��6�^��ٌ�Wrl���Mjl����l�!ō�Ib����o�D�'-5���V��t�{���1�����I�o<��ξ�M��G��RX��b���Z}������~��0�Z�uk��k�x����?�h1a��5��$N#�S��x��蚯+��/�m��|<EH������I
����C�� ��Pz��Z�Z�c���c:�Q�U�e[�4��4�XlxVHYEB     400     160{o���ٿ�    *C4N�)R���4 A�w*Ϧ��;,��Ot<^��Z�-s��БH��b/׆q��$�:J��@!��m�z��ʹ~P�|m��5�-�r6�XZ�Q��Ci�P���Ҭ�-�i�?2����x������Հ�Yk-����"��zWO����!WӪ�#[���?�,�x�a��W�aPS!���U���ܽbl�\+qS�f��J�vc��?>��(;����%Q���L�S�E[;���V�J4��O��4:[2�>s��:t���w]�B�i����*���ܭ Qn궅mk��K?r5�y��1f+(��pOK[vH��i���&���$B���q~��XlxVHYEB     400     180�6 �u]^��үJ����x���7�RH��5'���o�y�M��&c�w�2T���B���rO`�[w�f�$�e�I�W@���
��_sv�_��G�V�w�:�ɴ���X���Y
F�ũ6\ʩ��>o��]Gh���֨#�r��%@�FS� �F)��W��^�>�|�i]�f[�d#�ۤ��o<Y�X�ȇ{��-T���%�D51e��v/F��&J���0`�H��Bb��]J�ח��Q�!kR+�V�T�@>99����g=TKIKP�ܩ�D�jV��k���v�(�    a���_���Ź:��Ԅ�5M�P�2�.�i�Ñt��j�Ė�q�9u���T,bZ�:�������[�?k�}y�<U(o� ��aG�Wv�lXlxVHYEB     400     170����Q��    �&���y�����1�ry.�r;�l�NM�z�ܙI�^M �H�U>DE�>��W�}��0h�.Z�͖a4�~��D��ll�Ju�3�i�I;/�a"6�TS�@��|KБ���ޡ]Z��@���(�&���H�y�:��;��;p�6�R��^������Ş�EI!wW��R,@w��y&Y�gݦ�ps]���pW���\p�MVvfn�^���H꺺�K�C �V�z�@���h�.�8����j���f��#�f�#S�(R�&��/�^Zu����`9�
Ϲ�<;���D�kͷ��J\���Y[u�⯦c�y$��'� �ac�$+zY�8��O�{�[2�B>�l�~�4��`s幐XlxVHYEB     400     190a�4�@V"r��4mxs�i��s�a�T�S�bB��y@6�ȟ~<%���:2�
Њ�ou2x;��4    {��M����Pǽ�\�����؅������5�+ƷlѮ�^g$jI9�C�����I����ft��B��\���X^��e���(6����Z۽^��2��sߚ�'!qU�����ڡ�Y�G���,*{#���֤��Cr�6c|�J�0�f�Wӕ�DD���-e��X���.��%祭Q.���L��B����/Z��jB�M��}9�5��t�6����O�*)eSt5�����g ����6��s�`f*'+L\fw��D��{m~��&�g\]%fHt틾���a�o�
?����ֿ�[�.1�U� �S�+J�3��Y�����XlxVHYEB     400     1d0�����Mj�գT�䴭sQ��+��e��f�9@ �سw-�
F/�Onm�;$6w�_��    =� �Y_�m�,ר"\s9�iƍ�Q�²gD6����´���KCL`,bP{�M�O-J咇��v�Ԍ�!�ݴ�o�Wc&�áCԚ,|ח|�x��¡r1hmp���j��94���HQ,N��o,4�qC8U���b�h���J�G]&�9&���@ܓ��oV�ϗ=˪6����$�1γz����n��B���<#��v?�uٍ�i^<��\q�U}*C��\�k传��}zWhf��(�b��h�H6��s��0k��6
�*�s�����Ѭ!׋���c���^f��5D42WK�����߶h[1
)�}U�#�]5����a;�Q���fZK��o�^�y��?�YS���bO#>��pf\�� �L�=bK�]ox/iL���*�<ɰ8t��R�ٱ�<7XlxVHYEB     400     110�T����׵��C�޳�"�h��M������`��Pc�77Z.�����!^x[�z:l�����l%�.�bd2"de�e���e 青Nq�W�c����.����k
^�?��m_1���#�:-y����ګ�'A"�+5��x�����8�z��,�������{���5���o~�VGu}����'�%VQ�l�jnp�^cK�C�G���l�����-9<��t�rDg"�]y�5���cT{��`m;���#*��XlxVHYEB     400     140&�d�#!����&J��hl�EPk����À�-eo����y�k�����w�5�o��*����4[j��]v5��;nK�o�e/O���m�
���\�B�P�3��X\����I���$Y��~��C���d��>�� &�����s�b'V�����S��)�P8G�D5������y
��,%O����P�·v����^��)I!.�06K��Ur�u��i*�����UϿtflS    L�w=��`0��9&YOu1YxIbW�=�8��[Uy �O�q�\�qZ�3vQ�:�g6UM "�]�zI�6����E��I�[��XlxVHYEB     400      c0J�P��:"�49�Cy���?j�-���D�{b�Ò�/�!�s��DfGb^��ۣ�{'l�?v x߫�2������?�]�e��e�໊9�.hzB?Ϊ��`�c*���ﱁ���4��\�0S�]�>H�j��d� �    I�=��c�zx��n�j{$?�n��i9���GV��1�1h��_�^ͱ���XlxVHYEB     400     120�B���ʚ~0e�2lQN�T�H쭖,e�����mP֭𶓊��9���&*�������`�mi/���
�����z�
�R��D͵ރ*F��YJ,�x��k�\о~n7�!�/�D�_�@ȵ��L�� +���_x��M[���!E�����?�h��#�J\�w&����2����9�*،�T*~Muf�xM�-��´E�ֲ��k�0��_m����9�Yx#;���a�_�%����ly���Ƃ�5x̽7��o��H�3c��u���G�
Ku��XlxVHYEB     400     130H���8A�d0����f�N���d2j�}��5��3�H)���ҋ���A��(S]��.�.x�(�E��!�P�H�e�
��OoEwe���_��"doJ�O�eE,qH����I&�=:ڦ_֬����P7��R�SD�b�h�C6�)>�j�P�$�Y�Հ~jV��Һ�!�"�}��D�W�:��[#3C����9�gh4-LԽO"C����s��w�n�D���r!�gؘ��;vz���'8��@���]�:߹��o�y�a#�    $�}�`����B5ARDEiZZ�%k���XlxVHYEB     400     120��7E��+P� ;�M5��{wԦfQ��(�*A:�� 1�C!S�ij"�Σ|Qj97��;�MW*�E�f���Dƌ�0��:䂋A=������G`�p�ndӾ�J�^���V�4���ZB��P��J�������%�f10:��|vHaW[\%cX0��h�<���d[�I�!~�7��:A��#��It���G#�J���C�#�ȫr�0l�-ț    ft��A��{V���7��V�3���p7k(M g��;�[�1����~l�;If/��>��f�X�XlxVHYEB     400      f0!�E�s�L�۳�6)���򁛎ع����G[��9���}d��
?��Nx�`��=�r�D36"A�Qg76�����9�8h@.?�]���^La�Sq����{G��Բ���n�m�D�S��M��5��5G�vm<F��"�����d�=��V�/�b��:�4s���U���]�v����������~!?8)4B�E�h��S��NF�3b)��$ڠwqn�vCm���K��:�������XlxVHYEB     400     190��Ã�u]WTL��0�!X~�'��&�KV�f��,�R�|<~�~�db�([�ea@O��9��a��n���3=�q�{��T�����;�LuC\��9�n��T�ј���R�v�#�Z�O1u�B��W    ����5J����T�����ET�Htq�����,    �o�O��C*y��i�m9�<o�M�#���휱Ҿ    Pߟ'�o�$M�sC�s� �S:�w����P2�K�3    ���"�8g�&�����cYĻ��s��Dw��hE�&��)�f����9�=�~�i&�F�;'EdÛ�>��`������KYfۉ�gK ED���l������'Ծ����=~�e�Ct���p=Sbm`��a$�|wp��`<�$����I�Q�`'7�B���XlxVHYEB     400     170J�ᄋ��[���h�����    :�e���<���1ph    ���Y1�p�N�'��ql��N8��~��0� �.�z#۞�>R;�NR>J,~a'�ɯ+7�n���A �I�-Є}�@�D��z2�+��A��R���#������h������%n+eh�>��Õ�I���y���'BLX#2aD)��
J>)ׁ���{�C ~Ӎ��(���$W�ft9������M5���(�A��C�i�C�{�!,(�G4ڳt�卼�P�����X    �%ssm[5D��N=�"mX�����I���ܶ���\f���%/tΕ*m&y��!�%��U4;��ka�����:?�\KIF!A��XlxVHYEB     400     150
���}wOE>S)��=M�n�e~�Z |ٵ��<:(�����غ6���ѐ�1\_���|�L� �Q    �M$bOi�4$�9�^    �K�әDP���$B���/���|���hr���,L){f�}����1�b>U�����c��Q��:�%A��K{����Fu�� �T����RB���:���p��I�|�a�N/�����̑�}��
�Y?�����j�N�l�hE�=����/C���h|�`gq!]=sm,D��FHd    ���뱅���ǹ<Ё<G� �<'�:Zi>�n���    �S���'F�c�\
�T�ҡr����x�eL�:�AsF���XlxVHYEB     400     1400���i�G�    ���r��
�#e��GW��� ����I�����ѥ��SS���n���o.E��cqplA�q,�^=<5��s���tD����X�J��P�\㏟h wV���:����5�;*�:�K-r�DW�M)�<Ƃ.�"p��Є�EL֛��E��_j�0ԚE�<�p�=�J¸�f�?~l1��b�E1�Q���-(��ģT��dgE!��"�}{��v��R��a��g�=U��yq6Uޙ�k�9��F-�[c<*i8���������7x�j����~���8��� f���Z�̀�����jt]�MXlxVHYEB     400     1509��[48�{����/.<�kua��`����.q.�ԭ$WD,��4>�+��    �^�f{�h��i%����P�L����-3�=?�������2}�K�M���k�j��*ݽ%��|5��m#�23�
V&�[2\����~럓�޿�L����Fr+~qS�D,Ì �cu:�!�Ρ
��\K�H��S�2-���u@�Q��
.:b��-�]��������A�N�Cq��#>�>�U]^$�����l�ۼQ9>��/p)��;�g�����yv��{���{L�!�3&7v"����p��B���� �I���~�5��ʦC8�kk:�SH��S)IXlxVHYEB     400     150J�.�D�ߗ)qq~g��_v���yJ����d��ZB�B��G�|ͪ�����~�yUޒE/���T���\z�khѴ��1��I`���`U�ͷ���0��+eW�rtd����'��]E�xV�.f��~�����t���
�a ��S�o�(8��53�u�EReq�^[���3��
Gk���m    �j��`�I���rIAe[ξ y��ҿ�=�l�Ù�Ȉ��u �`4��N�W���D�)�(ΖU�[;vR�Y~��� � �u�6�yj'T���g��I�|�K?z�'U�0`�/�锊*J��
ӈĥ���co�F����\�5���b��Z�Yq<�/    �g��k�K���XlxVHYEB     400     130������Y��]W�pF~]����}��G� ��I��F�*��N�U��J���±�=��5
0�M�=d`N"*�I���]�tF���ׅ�f�D����^kF��z=i�|q�:�wK%��y=��%���D�M�D`0�Or�    ��!��:�����"m8*���<���3�����%���wW�N9�-���c�Emv~�:`����1T��E~�Z��L#xf�{M�=@�A���֑��� ��s��8���#B�՞[F�$t�re1nk����&�_��=Y���5f6�Ui)�q=XlxVHYEB     400     130)h�hDNQ��2�ٻ��m}�a.OGU�ݕ�45J���:{��L����O�-@T����Gx޲<�$�[��Fd��FJ��s{�sM�tw��H�z�7��U;��=�R�3�Ú-��K�\��Ҽ���x�{�T�q(_��_�{[:Iz_놮>�gI��w:ճN�ɷ��e)���³�����\V�sA+R@�ޯ��)b0Z��4C�=��,�Hmٸ��W���tv`!��D�b����A���[����7��g����A�l5�*Ix�B�����w\CМL��6�k�QS���R�>L��&(XlxVHYEB     400     130 2Hc�Ҩ�_Ąs������L�c�]{#���ڃ��!�x�+�+>�5����.�x���{*�7�q^Ԍ4�����>��}ϰ��h4�DJ��w{����|��R�#��3<_�I��u��/N����"����)����D;M    �ج�}-�&\�Y�#L헅6hGJ�;�h��Q/��,-�0A�c�s�o�M�T�G�8I�ރ*����)�h|�1    Z����<��
�o�g!�*\j4�!J�h���|�I'M�3&g���(��UWy�vJ<h�]
��k��Ä�^�/St��6�XlxVHYEB     400     100�Z/�B�sq��5��<��]\ʺ�C�ɥiM]2�0!�%�Z��^��������j�/ B?*�׀    AL��֖mE�Ӫ��U�h��*���{ͣr��M���������� �3�;du���[�����|����ˣ}�Qa40l�st�{p�p� ��&��n��y�|���2wo}eǼ}k���RId#m-*%��i����)hk�tB�Vf萰�#���g-�u/�9�$V�������H]0�+�+p넆���pwP�XlxVHYEB     400     160> �Q�}o1��Z��    زT����f��Ď���B��*� �d�=��bDx6o�v�rP��L��?+E��A�0�53�"߶I��#���D���������f|4�y�g�@��U�t��׽�ti�E��O�c�@#�ש[Z�b����6��p��-��N�8ꄨ^��V[ͭ��زo�v����Bw�ޝ��֌vuػK�u�.�9���h�.�����8�ȕI+�����B���W�2���3;W7�?E�(�'�ow�n��������h���#F4�pYzI�ۣ4U����S�7�[kk�[ϋmV��J3azri8��E
>E�i�i56�eØk�yx�XlxVHYEB     400      f0��S{��1�� ��8�����ŏ����pr{D���]6�]��2���3@_����K}�b�鲽]F4����w�2����ֵ֙`����נ�٩�=�GD�n�$3� �� ͗��,:�K�����<���$igpN�����!����w���镗�y�Q��MN�kE�ʇt6� ��Av���uU%��y��Z��/*�A��gl��mC�j(q���v%���o�1ya�xXlxVHYEB     400     1700|�J@o�.ɫ    Q}�齥\q*C��j����?wi��4c���mpq�V���� u�    �uyO��η�խ{��}������p�@�.�K���Il���������޻<�n���x�     Z'�t��(�S�����,T���.����,�VA��\"v���aSt�r�wT�'�~���)h}W�#E?M�8�1��z�AY����񋚮^x�bV�F9�`�?'s����.xۉ���Y�Z4�����}jc�Ug��j��e��ʃ8e��P�]w�0�D�>�|{M�y�c�AN|56/�����������/6�<4�i]�~u`*�=z_k?���}���CS~��H��CQ��XlxVHYEB     400     1a0HΌ}�0�$N��zE��]��B�뫆��hW���,c���:���N�:&��x��#�<�|4`�xEy��S���i��\�;Z�g�PU�#*�.߰/����`b�#i���YM�s����N�������Vӥn�z�38��p    @|݅���h�5��+    ����P�q�1�m�U������    ��s*"�ܤA[F��Gd�[�zZk�<����?���܎H]�W,8w����"=�~didSm�9�� �n�~$+�14��98��PZĹn׼m�j�9�u�6�팞0+����fZy(�\�KB���h^�5E�h�lT�-�-���ݞZU8W4D�@W�A���Q��ŴbԱ��%����Z��;M�i�o�Q���Q�    b�6}5�%�NK�/�r*�AAXlxVHYEB     400     1903R�B<wgs����;�e\}?���<�_�������]�!V �D��<�Ts!nɶ'��LEқk]ZɾW�[f,��qi��3Ϟ��AR���Z7BCr:1�~m�"���pE���    sd�    ��q��:���d�r�����    Yy�u�l�ܭ( ������4,`h��vY�(�:�i�A�H�à�]=�Q:�;�|I���+Vz�zGyP�5��:��!���?$p�s"��[u��Wv��O��NҺE�M��$���gB�f������R��`$����1��.n��    @    �ѱQkEBD��>u�����& ~D��a�A�Z�    ��Qw*xr���b��l����u�&��N�Ǩ�~������Q�L�T�i��%�^vwg�!�x�A�B���XlxVHYEB     400     1b0�t�N��Ɉ�=�������o}:?acnjN6�:��h���`��,;E�a�W�!�.�tC��{d��6�Ц��à�/�q΅ѵɫ������T
�q�a4��:\&'I�<��5;7߽"E�h���=��]>̆�%���z:�hX����(�>�^������&H�P��x��!~�X�����?�Ra�UE�YnWj�2�S��M9��W�v&�$�C���$��Z��Bax�O_B���J�b+�O����s�y
�T1�ڪ5�/�2iэ� TBQߨѱ�����v�"j��)LD���E�\q���-�a++w���j9�R�x#����]��.W'�}����WX�c�뤗��T�:�.����cdX�)�?{$��/� :�k#�;�������4�&O1��Q��)�����l�k��`kFXlxVHYEB     400     150M$���V6?X���\���vĔAS�l^1��ܨ�Ѓ��    {>��H�:aH�`���~$���*/��i&�/C
�fQ+>�s���c�����D��ǔT��K�/<rÆ�P����C�{
�z��FQr��L��:��f����d��z]����s#m��z�l��Û�����G��e̓��P���:�����Hk�K�!t�����%Y�V?s�"�    �9=��C$��v3L����l�Zb��(L�����+9k���7��%#��"��}���sf�!Ɲ�ᇒ��Xb=�(�x�Hy�2aUq͡}Z�->��L�~� ��������}��oZ�1���XlxVHYEB     400      e0o�~V� �b����L����>h�i>=�G�����3�:�g���ͽҶѦ���w�8�����^1X(v���S�4h��HC�ɔ��(
Z�D��g��Ԫ�!�v7��#����T���q�=�L���9�1F�����Y�$��.}�    ���@y�:�����!_Y�-69>��7n0-:W�����%�vqH�+���,@9܋�Q}1���i�]���\U��R�ʸ\
XlxVHYEB     400      b0wG�ڍV��C�!�^ȳ��
����ś?�a�T�<�7��2�'~�'��혝��{^v�*�2��
�&�#�n8(ي��#��"�L��E|��$�oƣ`��\6����L5�g���a^��ˆ��w�J�^�-Yk�<˽z4�d�S�jivu���خ��u��&�����6�XlxVHYEB     400     120�0K���`�(��۹pS���b ��ʪ`�q\����oȐD��&}�r�:,P�q{WSG�y�BrQT�QRkMjDVE�5As�    ����ֱ%U�[�#[&|�r�ШyS��`�z(��8���2��g��>�Ը��]~�m�T�Y<��`8￦�&�jXv�F�����z�b�0+�kP}�ڏ��$e���C�B�3�cч�Aq�J��<�m)]��H@7���˯�g���7Rf���?R[�ޤ�Q���Ǐk�>Z��.ڠ5��y�[�"�ـ��=�7CQ]XlxVHYEB     400     160�In�<=C��A�    Z�4H�<�%'�{0��Sφ�
&��n�Smz�}���V2�1�PE��Ty�剻�,$LH}L���陦������<�(��rT��#�F�
?�EĮ��-Tm.M����W
���+    +�Qa�x��07�ҕ����Z�&_��G�I��\��=���Z����6c�M�؁��⻅V��i��z�nI�u~-�2�5y�{�?��rHq�S#���
����q����B@��]�RĻ
��}��������"Z[DF�D���}��T��{��݁�r�j o$5O!�Q�U+2 W�̎�GM��m�ɂ�R�e���r
��˴���X��dϭ���XlxVHYEB     400     160��%Ae��VE������<=�ꎽ��;��-,��iY��ׁ��)��k�:o��e��7X��?��!tB4��S����Zl�ӟ�o���Յ���?$�^A�_e�`�������?9^
>�7{�R�/}Q�|N���4>A��7
=J��n�%���t�k%qZ�_��Z WT���w�]s��jshK)�R*�{�:6����O%��بj�
Mp��ƌO�s�>��4�[�Cܐ��˕�7��O�j�
�i�軜mL=�@���^_D�FO ��WO/����4��L�R�7��uH_G�2)b��e�N�o;Ԝ�SUdV"�8�9*��#0��b�[V05}BJ�XlxVHYEB     400     180{�( #G�6E�u�Q��o�[k�=��;���Jzq:���+Q����$U���    �8�;k���']�M�#�E��GcGXu��Q�v�xWC0d�^�*wv0�-R�\!�U0��e����9�%)6�%(��)a���2�Q�y���!����GMt�
>��j?Q�`���B�z}E;�{�U�̝��M��ʘ�zb��ۏ�P�'���=L�R2V�֌ST�������}H|v��;�����74Mߕ�ʈN�p`Nua2r����{��J��v��y���T�R_>bzY4�cY�*�X�
���j��/:W�D���pmٍ�rܯ^jH>��;��Z�q��� ���V���{vH����>�rM�����u��K�LXlxVHYEB     400     190p�7|1-��Y�����,�3u�a%z�x�/�lOR�<')����9�������p8��5��oe_M���|6��z����leAI*PL�vh��"w!H�Xb�q����yH�^=j���&;ջ]�wԈ�W!�.F������D�0��Kѱ"��[��5G7 �h�D�d�lT�2��9��/�r��*Ŭ7i2����$�6}�Ж����^�.��.+8� �P}�(@*)�f�Ǒ�������d'W2�<@1[f:�1_Q�T���q�]���0�th�A��s��    �([xL*1��
��>����2��e�LU���8����s;U귿�F�i�
��#C����5Fn�Bm�/�T#�"�j��أ�_�t�hE�ʍk�<��Z^D\7��mXlxVHYEB     400     1a0D��v�` �L����r�Wi�H�l��!|�`�8�"G\m��iQW��L���|���Z].���*�Y4P� "�Ը�ڟ����S"��ɭ��rN�q(ݦ�M�\�FI.�ޔS�C{��:"r�Լ���[��"g=5d    �ps��`H�_S�&��)i���ԯ��EU�9��n�F*��8Q����.��}�\��Wg��f��    &V�� A/
?��g���K}i"�4���a��d�!<s���<�cY�Q,�=f��$7�
|
�a�t@z9��ݓ2R�k[�ZӞ�<�ο90�>)JoJ�,����dfYއ��a�p�3����]@�4��L�w���s���� �n��i��Vw2�O�|�Φ���p�ȌҒ�H��)U��� ��W�
��Z��XlxVHYEB     400     140��zd��OR�Q(Y��8�^��}�V@C��o&J�&�ťJ9"6��U0mJ�Ln��fi�Nt��,!�����Y`@�����1��,���@���w.�Lڛ����&^� ��{Q�il�?�N'���O�m-Ƒ� a��Z�^�� W�i)2L�Dnēz�&����u5��rƝ���D[K�ZRE-b]B�\�5� ��L�V^F^�;�'a�佺K�2�.���Q�ԖR���z�0Bij���n%4+8g��27�[��o/39Ly��Ǿ����NZYpuU�¸9�|%L��Fn/�96R4SoT<�XlxVHYEB     400     1c0��ķ@B̺�`?��o�@w�'�[�JL�)�%�z��6��;&}�u�+�%]�y�Kۃ�[�ԟ9,����%��ZO���]�Y��۴�15F�R1f�+|�����޶�����o�C��J��?>�ϙ�Q�B�Ҹ�O���AK#�f|,�Ҫ��t�'<�1)x;fzK���o    �C:�����=W���l����SSG��l�}3�^DS�X����0�$�/h�u�A�窼��U�k��Si�qG�!�RMG�v��8�k� P��9 �*�G���A�l�S]��D�@�v�o�ӁWbG�i���Ղ���jy��{�
���,s�j�."�?��h����,C%�qS,$���V
 ���bz>���s='�h`w�����s���|\Z6�,9�$�N=O����Z`����)7�    ���M?J�=צU��
šz�XlxVHYEB     400     190,dv�%���́�wj�&X��W�8���,K��Xk�������/�U�^�,�֏0_G�Y����i�Yq�[��L�2��nui�o��8�yǇ��PP��s�S��H�Vc�!��bP�#�4qY��"Ƥ�    �����ٳ�ʳ��Y.66�)�ZRO�n[�˸�$2j��\� s���@�5��������S��������Bq&~�}
��-und�V���:;�����_�qs'��6�/�T�o�����hM� ���i*[΂��r�?�y�'.��
���a�q�;$�,X�H2����\D��d�,����F��<������v T�7$�G��ԅN�u-��ZD3qh5��K����?K�('*���� �.����Ԇ�c���XlxVHYEB     400     180�؇qU1]�L��u���N����������r|�}6� ��s�M��Ƕ�tZ�����e�D��e(�x��g�>��b|�6x0�;ߝ�������W�1XJ�gD��Ū�XU�:B�2��\c�����Ͻ�ʰ������P
������"=�_ �'޷��a������#���A�}��=����'9�0�1�5����5�5��K���)�o���Jd�J��x    �P($��]��+�ʾ�\��ye`��C�1����bx� �Qq���VxQ���z�p�^�9C�� vW�TSؾuiS    ܃�">t�"'�hٱ�4gK��|�[����i�U���9�yBm�V�����<��%��*��
P�?�0l�1�XlxVHYEB     400     170�v�/ �'�3�r�]|KϘ �9/f���(L\���@��*����$���8w���F}{E�=�c,%����\��G%��w=U��x�X�)�!����W}A�@��7��������!�f3:���!!J//�H����ԗ}��Au©RaW�F<6�Ue���?���<�gґFey{A�l��ɥFS��l������t�A`����ك�����Q~���s0v���j��+<�n^�    �Y����D˞3|q��l���)c��BnIPqK�(�/R��v��N$ؗ�+
�    C�a�D�H������g�t�0P����a��(��(����pǕ��p˒�8L����Ě�{x�F̾[X�]�A�XlxVHYEB     400     180Jij�9�Y l:����L�h!΂����{ә`�0��tZ~i�����e���s�:%�0��\㚅�*%�CǬ)�bڕ9e�SsɮL�@���9#��m()��p��:��?�
�$zhe�«�~�|r)N���6��Bh]�%ɯ�ǅ�p���ZlzͲy!Ї�zqܰ�����v��ɮ5�-�����x�E�[�<,�c�����T^Pܶ1Z"?�*�bj}B����չN��I��w�>kp�ܵ'���ɓ���t�"nT�tV?~��A��nTB��X��-�V��+�ԏ�-����uo^��^��b/E�����c���r�����S��_��G��Y�dN\��,A&�PB5�����pf&�]�??��Y1�jXlxVHYEB     400     140Hm��9��v���7�ZD{w6����+uǹc_q�V$ ��`� �L�X� F,�:}�`zj�#�bs���v�#���|�/I�j��d�R�E�s�_@�0n����є���\���:�    ��K�Ƹ�'\�:�l�����Az��U�g)�1Ip�ۊ��}��v�q���mu��,��%�����F�j��w��5��qU'z��>�>�m��6/a`q7�1���$[�a�ˀ�t�?�r)�u���ӹ���?��Fa�Y�$�G1u���;řop�~ȝ�~U<���֟��_%���b��� ��25w����.o���Ҷ�XlxVHYEB     400     170�&xavCZ���B95�����fY-��'�Yu��T�(�30Ӧ��\�]�����&q,ԉ��j�i�ѡ��^>Y^;ȸ+p���j�T�N���k4��C={J��vn^����mT]\������Z$�i9� \�{E�6صF�[�>��מ��TcH.itފ�
��C��Y�|a�A!�`+w��.J��O�g.~g��+�@7�E�Se�W�ܰ�슉ĩ��1�
���X�zD�q*#u2m��s�fE��_>��'�|Y�|�&5YI�E�j�n���v�)K�a��v="�3��wQ�L�V8��Xh����S��u���Ef��\:|�D�_$-Ӹ�р��%�$m�Q���u:���t,�l��
Ƙ��Q��YM'XlxVHYEB     400     1a00/��ʌ���$�n���)��sr����Ң৖X�5!M{F���Cč�[WҌ�jK���j!��1���9��d�
r&3��a���_��F��J$���,��-Yd��`�����܎I�V}�@�|�C���2A*[Пg�i
}21��b�H    ���H��x�E��ɋIZ�3�q�~������Jb��F�."
�M�i/z�)�]!ş{M�{;I�E��bX~�������U7"�m�V�9�p?�R��S�D��3@!v�R�#�Δ�A���Q�w6�4ЬY��*���Q\h��Ny����XÔ:B2^�!C�<gɮ�;v-׾�    �v�xl�k�/G�aR�q��sƦ�{��\��3�\��L̐$��e����'U�賐Ls��h���׼k8b�S�%�S�(j�-d�UXlxVHYEB     400     110ZP�#(ChmK~/�J �����@1��3y�(H��HV�.��K��c�䭎���{D���[� ?�[~ٙ���o,F|��6��(������2 'YvpQ땁uܑ��h03�Ktǲ,��'���'�~z~O��+M���ˤ�R�m�$�J7dCy�Ǻfi����A.hG4��� f�hĶ��YT�|�锷���;6�˷k�,I5����wH4� ���p�m��`�tk���Q�&��nZ\)"(xQw�^��!�    w��<ba�s2XlxVHYEB     400      f0%U@�n
gI׬�6~,z����� ?ϳoQ��G�
� (j���jJQ��
�Y�<���$l��E����J�E)�|J����!���`7j�*�=�f_���]V����SS��g��B�uNW��K;�Ǆ�HbMZ�i�2�&�+H�uh}�q1�� �Љ7$_�
k���#�kԛ.�b`6`����J�����/���wX0�
8��n�?K"�G��9J�]�m塧Q�Gke��y���XlxVHYEB     400      a0���E�#f�������J�k����ݳ�7��j��`�6� k,(ce&���]=I��uX��^Gy���H��>����|B��rΒT���px���`9ԅZ�B���q�� �&ƫO ��*w0O��KsAp��4�Bs����y��1���XlxVHYEB     400      a0��6*�-Y�c�ܤ��?�K    [syH��ӱX������d:���<�!���'��CEDPL8rw�-�g�Ro%#����bS���%!�������џz�G�b2�v�d��r�v�~5jeC���(݊ǈ��7��4����M0%ݽs޸�;���    ���QXlxVHYEB     400      d0mTSPE)�/�P%Re���k�ͅ
?u�I� �b;�Sv��1�ܛ��6_.���l׭`�YUz�u�
'C��u������d�&Z�\����;�H���G^ވ�9�5"o^7�{�޵�-�Aѻ�W�n;Sc,�����
 �wJ�3R�dF��ʬ��{�ހ�}����!%s�[?R(����i'�:��Q�뭣��]��#�jhhH�XlxVHYEB     400      b0��������FЛ���G��1_    v~�#��ŏv~v�tVQF�|J�/�S2K�n�dH�&�Z �"�����iǐ��    ��x�\# �0l�b��5����}�������:a�*�\|����MhCw*���ã�4o�y�n��!e�j?���<��-I�u[5����P��XlxVHYEB     400     140U7�]�.�4��;�.���7!9���@!w�c�s�C,(��<�I�GC"I�^w�É�nX�t�%(p|\l=\ͩ�0��!9@�g!է[��0"3��4���B�5�j�c!�wZC����%[>�ĵ�}>    l �M�ݴ`#�+�Zu��WH썈�8������@�R�"����dу΃�=ݚ����)��~����L����`�9J��}_�����fW<���ize��5�
&��JRୋ��QI�����wu�X~Ae�U3qV�K���P�ci����j�/Ճ���q�Q�Tn�?�G<(��"��ĢIUXlxVHYEB     400     150h�\c+wH#����F� �^^�TT���=]�Y�u��QK=�&�6h�����3��7t�DyW����~���u���s���7�̣`�:���Ώ���z�0LR�XQ�)h���&#-I��:H��WDb7����GB�P������F�`,�Q��͊R���D�����+h50ͺw�q���{�Z,.�F�r��N�)��?7Z �n�>��c?3̕���/W�UZ��;�i #�6��'0� zD ��|\б��܄�,��N� ��x�}��J�:����T
���c|��ᬜea!��QΕ$4"�'n���}�j����{�[+7�d�g���ߤ&��XlxVHYEB     400     140�om�fl�i�_�@���>`�i����)[~C���#��^i��ym��"�0O�@Jg9�:�˪7-�^@�f6    ��sN�-�����������<qU7����!R�ޖ�y��rμɏ)L�b��(�oG\3�uM�.Ԑ��Ȉg�o���:E6�`�:θ]F�Ϊ�.��=y@ܳ�Y�WX �4��P��SJ�s#^u��[~�XZ��������M�6pk�串-Xond�GCL�:C��
.��V���-_d�_|ua`��}�>ea&^L�W������M�oL���1@R[��M�Y;��[�v�XlxVHYEB     400     130s�3�T�/~bO��:�4����7yD��ź����'p��c�ҩ.��Z�WB&@B�
!'�^p�0�X�$��0��v�y�K�����A#���=rf/�F��k$
{YOd�>��.�6���ѵ�g�Ɏ<�ɀ�I&\LZ�)MLautA��ϟ��b�!KQ��ct�2̽V�(+{��67�M��͟ʩ p��p�ө�ɲdz���
.���Q�M�a���g{3�a
�/�풵L��h�y�"���Axj@�e�~Q���VM=�a2���� Ţ4wo���EK3�-���(d/��;�XlxVHYEB     400     1405T^�3�6��<�MD�J��٪y�R(�f��}�G�!���c��M�l����HB�R����FR�,D�.M� �go0s.��d��3�" ��솥��J�dE�D�邊-p��z����X7�G��b�*���b��9W]�r;�@M    t���nǯā$�8y�E�kA��te�(&xh��b�=fAB՜�=�� �Ss�����!���$�����~���Zv�$|�M�u; p
RƩq_y9M^������a�@�²F&*����� �s���W�����t��x��l8Pq&�I��&�9�m~�7��x�XlxVHYEB     400     100�9�$��<����n����g����'��깲�^����Wf��ׁ��ىhZ(!1ߐI%�5�b n�9�03�v��2 f0�r'hNn�W��~���`�mE���|j�U&�#�����ϭø�8 �������&�l˖n��ť����|}������p���ѩnM�_q��@f��py�3��X?.� ���M�R{*_m�:�O����\�iX�%��TsZv�GˎF���2�7Q�TpA�W���l�\ҢcA�XlxVHYEB     400     190N�xqbd:Gy��(�H��F���M�>gn{��уԪ����̛I}������J�y���"�Y`��9aI�n�LUj�!��4p�J; �(��/���;�t�XE"�`������D��ꏒ�v��
`�]�[�=��W�L�c���R3���6���8�z%�`�?���2��ڨ-�z�:+�~��k��$�O�)��e��*/��>��S�b�I��7ߥ6�Em����JI)ݣT� �y^�9�͈�1X7�\lsPF�<hf1M]cq�-�����P����0�y�Y���:�ܫU憀c_R���2�M�C� n⻘�&=��p3>�iqjɋO��:�������g�)    ��f����x�h���ȼ}��'�(| Lgb�����zǾ��@7��c�XlxVHYEB     400     140_�q�A�����-�극�b�VG�+�`�F��������������?\B�yS:b�׾j�M��J���d�k�ẫ��e��
߆�1]g��h�҅I7P2@�,U�JȢ�+��3�Z    �ERf�C�Oզ��v߼��N�$2(�( �D�(��2y��(XbE�r�S�� �ri��t������,%���Y.�!%�U�a�V���C@�W6�9��;�?=�a�;7Y"yU|�����r�2R�q(�'h����C�.�<�(�:�aΘ�$n��W�mQ5����k����]�5`�>}������4���������9��XlxVHYEB     400     130�`XmZ�a��q���zUr����*��[sZ֔/J�x*�a����ׁٺ"ش.��\�e�#��."����(^�̸��    ���C�}����m��1�q�c�H]-I�!��*��Tמ�XҮ�Q#��?-��?R�`"�(�:n�UL�Ts�i�F�����.]B�֓\���3�W��%z-g<�R�.���w��% YA���6��V��ʼ    ����fC�M�w�}�t��wR|��#��Ȭ��|�ʲ)����3M$��    ��N}�ۅfO�X�9|�o���]7�:���s�t�1�XlxVHYEB     400     140D^V.gzCƛ��8��]�a�FqW�>a��nP�.�A8bQ�ｎYM�~"jҲ��r��q:L���A� &�o�7�����    ���79#m n����t���y��AK�{/�͌ق{��L�ܥ��80�K.@��������ט!�zV�� �r��x� �ѵ<��f�­t_ѐ�H~,e��< ���y� �9dx!@�    ����#�����Ϣ;Q~���̀6���GRU3D/$�|`N%�|F�Y�r%V�{�'�L����=p�O �'�N~����m�[�~)�Hw�L��op���z�0\M|9��h�XlxVHYEB     400     130��XK$�X2�$O��)��bO�5��"X{�lA/(�oޏi��35����h���i     �'=>[��f.��B-g�����ϫ�D���Er}�5<8@Ȳ���!V��l�.�͂��䚕4����:��� ���|էc���k���Xq�aЎ6��,S�?�˄���z��C������zS_�j��&���ŕI6�y�!���������|�k�x�mt���J����T�}�|���i��YXaY���+���n��t'!U�7��h���Jz,^�7B�v*p���-�+���5?"�KXlxVHYEB     400     170    P[�M�;C�~�F�����vG���C��B���G(��*���OC�i���f\л1�hC�gR4���i�OEp~�    ȼ����M�u�1.�}u��g�r�1u���`�    �S�@/%��NB4p��ſ�����`�.�y�F���܊��'�s�@�P�$���(0��Ӂ{�W��1�I=K��b���Ɛ�W~�g�6��8��,|x�vC_���    qf<SN4������ t_ !*�?�X�|���`�No>�o �B3M-��'�պ��W]I����[��|����p�S��Jկ����-�1����<�g�����JII|��{_��lc��nQ��M�H�Xp�E:"�:&�\hXlxVHYEB     400      c0E��7]��d�eÁ    �Z�o�    ���f�����goc�5���i;S���H�:�S�쾫�_�*n�{:O��������O.�}G��qqDvs���۽T��3ٻa?z�
�Z��VY�ɮ5/��vmnؠ��ϟ�*,WLy�Oz�NV�3K&����#UOD+>��lL��D.��m���7-�oRXlxVHYEB     400     170�V�p`kA�B�/t{� |��oNƈvb��m"��lH���,*!F��`r�ِ��?���=�"���+��?Ռ��X�\��>    5,����H��M5ڸ}�c����_<l3h��ge��"���v֦'�,�$Q�d�9 f���(,�a�Т�]H�J�i��'6��4��~�S�m�u��m��l�߶m�U��A�] ��]�%ݭ��S)�j*�zC�d��x
�ɏ^����fX��!�=���M:�;��e�4�b���RH�p�K�z�;r9����e6��ؾ�4�$\�t��?��J�Ӱ�C�'�Bf�!(4�idh!됄��B���B���;>�My|봧v9~��-
�l��RYy���)XlxVHYEB     400     1907�cͱmC��+��+�,?���W�0Z�����G=Cm��7T��΅z@� 
�3�
��$�8�_�\�˖V!��<���R&>GA��#��O�J����R    :l���x���?Q�Q,9b�(�l:��ױ�eO'�P_���P���B��m��pqX\s�ű�+�WD��{.u���W� �E�?�����S���K��Īɴ5IG��#����V!@"?�_
�F���
o��@�ho��<bng#_�3*U�/�MU+X*l!���<��LI��3ńM��S�}+�S��h�͢I�S9h���P�d�p������fCN���/���?���y�� �`]��:��S�I�H�c,�:�/�t���j��/z�vX�L�Ȋ�-(    ���*��:XlxVHYEB     400     150���zy]�IL)Q>��͒��t�e�n�
#�-��v=:�'m���W�z���L���cԕ�V�K�Y?B��G}u>�P̝�Y�;+ga���J!eK�N�Y�ʨ���a0S~�͗�׾�3Lvu�?����{L�5ۧ<���W[r��[��ڃ�=�%�(��A+b�lRA'�)�.�ΐ�3�Y��H51T�9�ܭ���a�+���m��B���U�9�Ҽ���&5���!�OC�G�Lq�3�\¦z}���A=�����L���|�    ?J�tI��,�    j��L�2���D���;-�
JN1�H�F�;y��M\���9�Ƴ����x^���XlxVHYEB     400     100%3O�x@�?l���q$��"�f��    ����:y#�m���u��F�d���٢k�k,�;e�,�bE�V�k�8�t���&���x)q�\��<��m����*w �Q)t���T-!�P�z�Э�i����Q�c8p��5YfE��Y��o�y�12%�+�CLy8A��~ ,�����s�q�P��_��j�L�I��d�a3y͕�Yے��'U`����c    �S9����~ 'E����^�m'�goa�l3M8!mZXlxVHYEB     400     120��y��m�W|�36�=P�lY@�����,~����(���)Uv��V���n5�H�pN��t`bb~�x T��6����0�Hi`}UOW��d+Ģ��f:��}�R��3���''��"��iK�{K�zt$ʻu��{����&���y.!�èqG�L�)����]E���@�lD�    뻪_��u���#z04�w�7���8ۅ0/��d��3P%� �3�C�n.��$E������[�!��}�.�~Y4tGVd��`��&f��#<&"��$�]MXlxVHYEB     400     1509l��־;�����Њ�W�{�)UM���RT� ��>��p�hxF�qu�5�@y<�28պ�esѾ���7X�
[�t}�������~N�wCL��}B;Zw*y��z�WcQ��>L�ӊ )P�)��2�a!u��>�6��0u�bޑFю���A�}�TK�&�8�"�����/U�ܱW�3�%�u��N���z6�p���,��6�Ex���3�vHql��C���D��cG'i�1��3_j�f,��C�k�Rt�e�.�Z)�@
��������I���JsRr����:��Cw�������=�����
O?��>͒@� �AXlxVHYEB     400     1a0&~�&l�W�?��qЅKU�E*��L�# x�H���NA�8���CY-�Do�Q�����uκ���\�$���om?9I�NG���]�p�� ��(��Qx����|��`L���Z��s?�=%
b�8b�΂n��51�!y�+�8����ɟ;�76b�i_�/��5�����mnB7�����7/�<mHn�tf],ڶ�UL�P���w�"�P�i�&�+*���k+�1a&M���`�m7��T�ЕUY���8�K��f�p�cS�"�a�KÏ򃛱ȴ�07O�1X����ߔo����h /9DS��P���)��t�4_���{�:FH�P��S/>�{Ą#q�)�M`����d����q��ϭ�q�&S+�eh�����4�CG�0M���o��j�euHd�CK���@���I>�tXlxVHYEB     400      c0Q櫫�_炖�`    ��b�ce���p5����K��)U���d�B$1�c�#&T00�Y����[h��-���%J8"���;M����eHP+�R��e㛶���3�RP(>m���ع�wQ��$Ό�u�u�\����32X���O�9RI�@�Iel��BdN?utN1F�=�޸    m(�i�����3��    �XlxVHYEB     400     130������r9���zE���y��E�e�E�`ur���VX�`�`��=FQm����0���ݞ��o�0I�J=�vV��SH���q���x+�+��\H��3�:F8ș�HR��B��̓�ND٘����<!J���bt�6a�<H���\��������Ǟ�2T���H����:Z&���8�3�GÂ;�{���i T�H!Yt�(Kzt�Q������͐�|]�y� ��oV#�肫�pCxEHK�vU-��a���N�۾v"�ܟ]0�җ^+�w��U�1����jQ�L<J�RU-�q�ǒXa%XlxVHYEB     400     19027\�(bـ��QR܁��W����R~��΅�Lg��6%��h�.7�0�    �����BEx�����C�|��3����ѫ�V}������/Y
��r!�mlr����w�K�6O����6B�1q�^�KT+�
��m?�N*[�S��
������g��mi�$Z^N�1���-SP�n-���&Am��{n@���Q�y�W2_�����=�'B��2;��G���t9E�Ú��ޭi9|%a�X��
�6 ��-1`˩g^�&�%���O�    #z�����O!&��ZZ<��_!��N$�H8+�^ήV��S�4��M����8׉_�3I$��bD��"�+ݤ��--�oh-��J�e���hQ�    �fO�d�$�<��:�j�oU�P���[&XlxVHYEB     400     190�}�vX�I�ÞR�j�����.�>�}�X��a�N��^�_瑧v��.%�}��!%�9�R�̬ܧVa���>��F�n�嗭�#X���6U3Q�4>�    ���!)��W����5D�.~�w�Ek�ݎg�õ�,;I��.���c���{:*    [��y�����z�T�D����Z��l����m)��}�ԝٯ����S��]�a�k�#H"�Ү�ܘ�ĪdN�7��W�N!�K/Ĕyы}l����#��*�$�
�t���C2��^c��Mu�G�\��.64�i�?֋6
Z �=�yj�j�~NN�3��?�@�
Fã�ޤ����+tC��I�4!�%iD"��6�_3�Aj�Xu�좄���?��6h̉�f�l��"�]C��#�x7XlxVHYEB     400     1507i� ��v����*!/j�l�����?��5DQ%@��8[�e@���d7�݋����쩧�&)�$���_²�ME����܎�:I�>C?yǷ_�P#^!�1�$v����H��e��s��u��H�����]�\���@�j�F�~��5[SS��,���op��`��=�{Sa�ܚ����I�;�����j�[ޤ ���<�B��[�&� �!�mI�{��z*г:� �!c�/[#2�_�U@c�u��_��4���f1j����{�<s�O�g��5u��Aj�l�h���A�su�Ƿ�07��t�T%�[�:�.6(2�D�0Y�<��XlxVHYEB     400     100���M�P�M��_3��$����/2Gx5:yZ��3�}5xS� �x��    ��m̘\8��䱷QN5;I&�E��L���82���ۀ)orO?�hZz��0�G{�k�K�\���9pu��UQ���Vkfz@���3�ߢ��Y�7/�����Ϟ�ۋ��nS�.���p��k�`���ҏ���@f��lz�r�=��b��{MU,���;���;�}�Ё�E�f�g6m�v��D�$��6S.�XlxVHYEB     400     140N^��Y���i�H���镟���w�x����l�p�ܪQ���P�$�:*N��y���O��L�C��gG^F8]�z�P�̮�?\MR����� �-�t�UBJ"|U"rХ�u�kr���6d�����w��v�9�����?�*Y��>L㩯�dT߹��8tK��?h�H� C���a�&Z�X`�\iB�N�3�I:���������)7���Q M��-9���E�l;�J%�;_⦡�u� �H��|�2��C5����gJ,�m6a:�2�W�Քn��\���K�TH`��Li�� ��@��d(|���%H�Kq�>�S�XlxVHYEB     400     170=��n5L�K�|IM���Y�@}�����M�o��M
�l����i D�޿�ֺ��w    �W_��@�M+ɤ�"���ւ�!{Ѧ���xu���9tX�Ep�iì1]�KG� �{_ͭs:��,"�Y�ZI�1D���H���On���iɟ`�Q�Gu餵��D�L�n�_��C�DV�i�ȭ��H����4+��[,`�d{#�ApUݥ<����l3Z��1"|'})��9$��s�p*ψ����y��6F��g`s�]��j�!un��v<�}���7�jg�)�#�Ö=�@���Q?v�6    �l�;= ��D�8V� �������SU1�!,w�EL�5�Ap�C���.{�18������ ����ΐjXlxVHYEB     400     180v�Uo�t(S�Z���l.�ؼD�/��jԣwջ�;�\�K;U1%p����6ɛ�Z=�����,��}�)
�0�7~wtG�����}\Y�Go�ӡ{��x�B�,��7�֤��X��hP���F��ǋY�6s󧍆���&����6'���X�t�A f��:+���J�ݑ޾1����:k��>��4��_�����F���Z�g;0���V�����������+>�?bn�hiVao��,�����F���T��F�ʃ��C��F��_\�7>
ˍ�7E}���T��� �}upZ��/R�T�ǎwR��> �rlލ�"�6=��N��u��p�؋�
nu�mC�r"\UX�I��Ƭqp��̐)EYAsa�{�XlxVHYEB     400     1b0�KU�E4
ٜ�/���;�������)��V)��N���XL�5H���fRB#�����-��6�L)���a����7J��9YH�܁.�y%���~��΂���O���Y}C��t@��z����jP��(x�ڿ#��'S��޶w8�3��JO2' �^���ңIX�{m�)�a��U�[�P����bw�h��w���Ɯ��j�^���M�����q�ROv�fs�Zl�    e�;Y$��6�6���l�S~`����O��HJ��zJH����%�*��y�5)��n �����f�x�㖼��S�K3���(�V��y��wH��"l��&k�`�a8�}tu*�s��N^>|��]=�(��f��b0FܪJ{�3#�b]��8if�Kb쨒������cň}N��^�K!T�,=�{w���e���j�忀���XlxVHYEB     400     180WTO�~    �G�2ݠ����[�):��A,VS����_���_W�F��M����M��ҮvT[����,�<���˅�7��nȐ�D ��ֹ���!��w��ϡ����z�BP�>`vN�i������
�,5�]�V+s�� ����(�����i*�IV�
����N&׺��{�����CO���&�h��P�W�Ϭ"��0Ws~\�    g�.�7Q �7}��1W�s!�=]v����UL��Q!]�f�Ty+������§���A$�7E?q�xu�� ��n��Nl³��lkN_��]�0���;LE���X@E���m%�^L�K�B%��9^Q>,����qS��^Y�l^ i�������c&A ��-|�It.�ll�XlxVHYEB     400     130�5�b:�cA������y���[՗�zKXs��0���>�_˩'�Cԙ�P\?�v�,�����F�}q����A��roXFB�    �Sd��e����
����)f    �ĩ���ssa��hy�Ik|U�>���j3����8��f�T#��'��B�o퐫���f��o�6@�B�V��w���    ݘ�[<���J��װ N��d    6�6^i�6�CZ��|     ���W�ۓ�~    :�]��9k�Xc��ɕ�0L��?�\�(��Փ�-�b�E"/�VS3��i����d(�������Z�h�U|+9lC8wk]�ٷXlxVHYEB     400      c0�Ie���sH��I�Xwd�\R��aˬd}0
գ��HOk�����{/�lM�Q1�l����
@ն���l�kgll"!���;�w�WO��h��WF�����b���
�v�G�(To����O��x4�O�ʭtG�m�2F��a�%q4��"W�*����g�����&ܬv�l<�x*XlxVHYEB     400      f0���I�/�>�|��=l�|�V:���X���C����_��f6{���o'�o������Q�4�<��砚��j�����_m#�D3x4�E�B����C���Xp_��ꟑ���_Ȫ��ɱ��Gڒ����h�g'5Z�
���t���}�uU��cv�FE    ��.y�^Q;���z<4�X�������6�|��ίn�.�_�d�C�D~i�    ;HQ������K(#/4m���XlxVHYEB     400     120ç{%�7bɽ�_&v��69�+),-�E�(�_e�.�/�~o����)DsD�Z)i�͕N��zdq��ݩHL�A�'��vne`}�9����v�����2I%-Ua;a�)�٥�z�['��B;�Sh,ZCH�h���޲�<��Ɏv�NJK:�e8���Q?�VF@;n��A[+e�0;������3���s��`����4�I)I�d�p�mĸ2E� ��&a��{b$Sz'V�Ń?��Ô`q���~a��%�E���p�q�6¼$�Ld�@%m:u�XlxVHYEB     400     110[�}��җ�.���3F&�D�F{�BD��cɹ��#H.n��w�!a+$o����m�n���*�e-F���+>��iV�ٗ��>�.VIk�f=��9\�����?�nV�    ��\Y����vxs?8��q��m��2Ɩ��|�<G�m�-{���E�+�+�    ������Ms�+���w��9{|��*�n��P E�6��[Q@�ː�Ao�#��HC���a|�z�������̔2�*d���j����er�y63'P�XlxVHYEB     400      d0+�F���]b�qTٮe)������PmF�[���.���0�˻�v-zm{4V�OJ{_��˾o�b^��d�\{���`� �g��Y͊V��@��x�i�\�z�g�_�,b��a����� Ekkg��8��f�ϪN�� �rn��SL��L����}F:9�"nM��؄���D{]`��?�y�5��0�2.�I��������F�ߨ��e���l!
�uXlxVHYEB     400     180p#��7�BJ$�ă�%��wB�G8{ C���U���-%�z}/�
m6�E}h/�˦j�s�`�Y<�u�``��)���ڔY�\��]N%���SdD�ͤB�� ���D�ћ�bt����
Yu}~��~�/�g�-<˘��������ղz��p)�����z��,�$��{�v4`��=���X(�+HIdvϠc��v�/�����ʚ��8�5�!j<���n�v��t^��p��M.�o��-��<�Ց�e;����9a͒X�c�>��׻d�b�����,�2�QDB&������O_���Ӛ��&�eO�]7@0j��5�cv~H�I�m�&J�F�J�,W�4[˨��;���{�ݷx$%�`�� ��j�B�{j���XlxVHYEB     400     150\(������0���u���-<�<<���?��PWLv�>���s���Ķ�"k�qmMw5i�bb& ���@U N������U5:����nf0l�ޗ�.�>��s�5��j�x���>}Us� ~RT����À�FE��� �    ���x�ݍg��Z�|4?��f��.���Oi�U���<��hw����׳�t��q��A������G�Y�S`�}lY@�?��P�qdC1��    �a� *x���n�j��>��Xx����|��C
�kxv\^�Փ    ȝ�����$,T�h%l��    <�0�E�z�H`�p(���7������lvh����XlxVHYEB     400     130p@]~:    ���΂�:�h\>DW�?�v�7����a�]����k���� �G(����8x�����Qa�\�N�G�P��~@,Ui����]i���)6����OϾ�����H=_���{u��*G�Qh�^�l؟��*֨dj�*5�U���ڣ4�d�F���9����IL��R7�#'
��F�X���߬�����\��(�䈞�h)B� �,�?�ٝ\d��ۈ�w�.��2H��r�:�.�*�r�����~m�a�����t� ��AvƷ�9�e���E9ZZ���XlxVHYEB     400     160@$�G��[؋��W�u<fʆ��b\�%�?�W��ޅ��O�hK�T��!����Tw���yU��E�U���E��n�b�Y��n����4
��8��N6HL���������)Z�u��l���&�����2㫼�����hN���DXCD?�����V�'j�Iy���ۀX��8ؐ���$zX���&Ó�e;���!q����/_��G��8E�|��,u/oBͮK�c9 ���C��w-��/�I�l%N��l�;�L+Nɐ��mUw� ���K$�o��"�����0S������.[$$�!����]5�o'�}���.\�@���$.�����*{��E"��t����XlxVHYEB     400     140b@HbO<�rX6���_0��Lwt��4�m#Jb�}����R�{Eȥ�v3�aw8�B+��p�����0NP-������f`���{���.l�`P��E*m�4P���g��H~���?��8`�Q)P@T@��ɹ����M�ӄn��XBՂz+:xd^_���31h�=�۽Ȣ(]�`��4���Uf,�����:i�vUx��M�Wv    ~9���7���'�X��L�8|���=���\g�ak�ε����K�<�b"���Y���B[�eg��V��(y5CuFa��T���/�@��玐d�?�+��A��Cޱp�XlxVHYEB     400      f0�{(,�������:=    ����}F�D��uP/����<�'�~�4b잻���^�U��ҔQ��~�T��'0#z������Nܕ�4�]:-d����z��>�����"���F
t��`��T[���8`G��Qa$��ÛC��#�q�/�]�h �s��U#;�Ͳt`(w]�ŀ�@�/Ѷ�J�    6��o�@$,T�?>{dj��l֜�Z�b�/��}�/�,�9~T����
�ṛK���$�XlxVHYEB     400      f0aIr��gp-:�E]{BW������i��������i�BS�4\E�_�������(�G;��Q���,L@�J��.�Cg��L�~w���3�)�(�w�n�Ġ�����%�U5�i�6�p4sո9�"ͅ�1�+�f�26X���#;t��ޒ�8W�����V��y�A'Jo�*cbx�;��h�ʑ��fj0Y��N�S$�0K;-\�m??�u� UU��lo�kw�9��u�XlxVHYEB     400      b0��j    �d��a2�����BFܤ`)��)���Z�3���g���-�'��.�R^���i;��~��)T媉D��Ϳ��WyT7r{�渜FΛ��(R+�A�g1�Ɠ�P���=�l���2�))`�0�1Ue"������lԽJA������ľ������=��5���&�BXlxVHYEB     400      a0��6*�-Y�c�ܤ��2��$'pi����F��OgN    PG˅N��������_N�H.��
f>�Wܓ�n|�����O��O�O�sHB���OL��@t-� j��k��,��4�_f�(    ~Q���v��q e2%��IJ,ל��wvG�鸤�>��'6h�XlxVHYEB     400      d0��w�#_%���#��[�38#z�R$��p�hW��VE,q��P/gi|ឦ�Kq��[����wzp��ah+*�ƀIXx������x�-s|o�(Y;��T9�XGJ���-�X�D`��S�`Bf��>c:�`���5\�ظ`a��W�������,�%�<�+ᬥq�dy\�J~�çl|�m��@��KÚ�P���W�_宑�XlxVHYEB     400      b0���:�ʦF��½@�f�I�#��1w���2Ig'�ri����O@��s��̨ h����#�|��jes��3�6kK�~�R4����F"3�0���դMf�G���L��{���}J�qU�R�d����b-u��    �|;)^ƝK�x����VH�d�Jj�l�@���ԓ���RmXlxVHYEB     400     110ܲ�6Y�iF��8#���5���P�I�iU��K-�4A��x�n���0HB�oB�$�Y�����/[��hJb�E�G��J�b�dW!�͇<(V�܈o��{�^u>T�N    ��X֍Ǌu'�(qC�nRuU��:�G17��dG�en,�ZP�jSj�    �j�tɉ�    �'7�FR]x�IL��R�U��߶�&It�t� �;�3�VjZ�����4�Z��Y���t������o�h8ſ�y�paM��q3U����b�`�����%��JN�b��XlxVHYEB     400     110Ƅ��MC��^�/�����!��
� �\�z��#������c�A��Q=�akc���j�n���h���Ĕ���=��t�֦ύ~fӀ96S �T���|qrb�Y)q�RuEș[�cdI�H��|b������*��y�"k4Z�6����%6�LKTƶ��D���t�����h�\�a����b,���ZF���    ��'�[�]N����]�@�za����i��0��1 Y�w��/�My�YN��H���j��PI���,�f�AXlxVHYEB     400     130@7��u����uQ��,�%�    :ݮu��'#! �꥾��&J������ �
U�8H{,�s0!E��wcK�f�:�H{ڃ�;�/����2P��g��ӧd��!�2Z�/���t>�X y�H�!A/ySr�y��(xڦ��k+���1\w���/�"to7�E~�[�{�|V�k��    K��N��ma� �zxE�44��P&�e����r��#N68�Αt9�Ɉ�(�" ��$p4��/:�"��;p��M��!����.��Hj�'V$���=h����?JPw��9�-�Ϟ��S��UȱXlxVHYEB     400     110��\^�x�2*��R�H䦗x~�ҡ�?��e:�^���1���݆�w���\^��Z���L�5�Lw"�<���(�����U�=��j�9 �1H�D�b�@(mrք{o�pn>��e���ޣ0 :b5���K������${��q��j(�a�܁�u{�T�^E!Po���C;�����cUy�;�]�Ap�������w��l%��
~O�_�ujGʗ��}    �E��#R�M��:�b��!D�!xO�XlxVHYEB     400     100$��iN4O���+9Ig;���<Ԭ�oA6�����iu���7�S���G^����i�[}-�ɽI�w�َ�뗹?ʊ�O���(��i�����[Y-d�!�g�#���d�4��ć��ä�����d�V��;ei���jb1l��D�W�X�}���F8��~���8vS�Z�I�˝� 0-5��%}�)��!9�A���Á4�C-r��W�l��@L(��P5�̘K��NKXJ�.(Zᯈ��vb&(q����|;XlxVHYEB     400      a0�f9Unt��:����V-���1<>Z�oy�J� ���9;�zV#�N��aH�    `OMk2��*Z>ҡl[�V'&�p�Q��@J��:�V�X��~`|�'|H�I�9�>�cɴ�u7#��AA��.t6l�=��+��a zU5զ����.�[��n*���yvXlxVHYEB     400      a0�:l��yM��V�ܥ`z�)�!���5��Ւ�OD��HWc�{��6�'�[v��f�}J!�]�/�߅�[?ҷ�3�a�#Hb�-p�XS����>�����z�ؕeR�݇�:��#������e���o.va���?܍'��Ic�K���{>kXlxVHYEB     400      e0X�û}3�P���ې�{�����C� �ǳ�~��Ž�Azk.uSg�"9�    ���Цݖ����Vrj�16
���E_h�?�9�U��y�/Ƀ���Ih�')
.���Y�v�m|�mS�y㴏���H_,��s��9��cc"� >�    Yu���.�5J�L�"��h�o!8�����$��3lI��� ��x z<��b�1(��XlxVHYEB     400      b0���"���)�H�Y�V�3���    �ϡ�Q�����-��P���|�[�_iW��x~�g���:t�{��2�R$�m�z�aMu>�D��57��0�B�t�𑲁�{���*Y5x*��<c@����n�٦�Ǖs,�[8,��ɡ���Z�9}1�-���2��}�9��������XlxVHYEB     400     110K�8rC��Z:��XW&&�>ݏj+Մ_�*��ar��*�%�56d8K�&��'��A������c��y��yD�g|ת�U��
��F���9����I�����$}����DϜ;&��`ٶ��唉Y�w���6��D ]؈|ؚ��4aW��y��@��*ϐ}FS؜�1w?���E|�X��|l=w��� ŵc�G�բ檆������Đf�[W�{��������ت$��E���'    �t��$��)�= ���(1Y6B�(����XlxVHYEB     400     100���½Ͱ,2��J�(�j��n����𮻤 �D ��T�K�:��Pi�g��V+��"�ybOq��pO���q=�}��~�˟E��fI��k���i>&���l�J�=V%;���hVO
惍��ѽ�^�N{M(�C
�N�����.Z�r�4L�nMة-��b��ĵXLK���J|8V��c�n�ѻ߲������L���F*��%�ԗJߴNxБf�k��d����v���&eQ)6��z��f�?��ZR���2p�XlxVHYEB     400     180z�h���~r�>����W1���K�iW~�����h�+Yi�%�v�����"�z�h��Cp!Kם-8�hW�9e\�YL�^&{�4����#D�i��^#!���+2�>�egg�bL �����_�E�|
�l��(��}�O�+m|`QF�Lg��`�v@�נ.��ݺ�w-���ݎ�}����O��`��α��    jM.a�4i>��yW�oG    r0�#Č��|�el�n6�w�J^�]���ӌ�Yu�N>pP�����l4#��ԍ�\GU��|�Fo�n�h��4���3&��.�M�^}�˖�!BO�ăg��W�C�9o�8 ��4���{6dr��dP#^TA�G2p�p��YpM��wIW�9�!����MR�XlxVHYEB     400     170Q;���8X��po`b��:���s���:�Th�_t�yN��FSV�T��@hr���Y$V�K��XʜA�&g�&t'��r��1��N�.4�UM-�JK�~�1���~5�I�`��#���-#�c|�y���8���whx�sL6����    �P�E�&+��ѝk�QeI�@�=˕�0=n:�*LuP��ҿ%�\�AZ�cF]�X������D�5є�k�]O���E��6�1���Q���&!�ۘ��c�l�\9���:.��;A�i������۠*��d���`�x)}�T�U5y���#�    ���E�*�gĎ��(�gL�Q�o��j!��n��k�o�{��$�^���֋���MZˮG�^�bXlxVHYEB     400     140x�8�"��wS~b��B��~G$>����,���pev1@s��f]! ��
�8֯�����H�j��۱��4�5;k����u4����`;:���?����<�maM�ߔo���� �l�٦��ܣ�5��J�UA��<9s'�
��u���A�w��ٟs<?i܊�Ha�c?�L
��+_���7���¡yψ]s]0c�����Σ�I"jtg�B�v�p1���K    ��L5I�#��9Z�1ZG�Ԅ�(�}�k��[X�9�
�t9B��D��D$U��Y)x����'V�Y܄�2_��)m����H[�mXlxVHYEB     400      e0d_�#��X���q�A���]�U��9��Ӹo��r'rm�,����<���O�aD[N�Er<ix��f�e8i*���5p�+�s��B�2�XU�=����} ����S�?uu��� �L� ԍ���D���D����[["&~��J�=��{j��~Ş������ܼ�gMǸ%�p����������V��)!_��f�&�8��ʡ:�ٗ�+`C�9�9J#܅%I�+���XlxVHYEB     400      f0�6�9wƥ�����:GPc���&c�T?�����;������^c3�/�A�F`L��&_g*���� K��Ǒ4l��ش��rM���h<��,�Mz�=g    ������5���{�    Tj�g��
�|\ΙI�@�
_-F1�rs��!��pje}�z>;��ڸ�]h�� �V���s�_���r���V�b�&P����O<�'$�1�m0g4��]�VLh�k`��B�&�ͻ�'��7�)aL��XlxVHYEB     400      e0͎�JGntE,Y�����n�2��t����wMg�����y�{�    2��BfvcO<M_�R�j�Hjn��8���D1m���3�W�1J�<0�1�˼�����&&��|��C������51%/V|�x7��*UH
s�r#9�_�U��d��wJn�"�6���������K�|�гPt%��*3fj��B�t���y�{t/��Gnq*��F�%B[m̢>��CɷXlxVHYEB     400     150�!��9���#�� �=P��a�N�Yk�u�|=Aa��j�/�ț5:I����@c�E<�����;��|�5�(e$B�K�
��锆W��b5t:q��2C��q��X��A������b7���"��U�P+�
_xM�1����Ah�0�睲�
6Z����Zi%�&���@��N��ѩ0��ͅ�#FW�IxC��q�|Ķr,�4�=⚒�[+V2�e1�r ���������Y�0ΟQ���t��]�'��^�v�%��Ng�l���)zi��dm_׫a�1�9��/9&��    8P�"����[��x�]}P�1x,���:{vX�1���XlxVHYEB     400     150�G��*�~��͛�(I?���ʓ���(�~�t�ٮ����!|tޛD?\R���DWc���j��K;���6��(&�9k��+[��8�)�+O
y�l�F#�3��\���G&R��'R����#���_��૦^�9b'z5Y��Ňh��i�ȣ\�!�au�?�h�L���!�A����
X@%BO��݋=���5n��*��/L]�+8����~Lvx\P>1ɻ@0o[�@
�Y��ۧUJ.���Ն��`�����v0'w?L�����u�G��+S۩.U�����H���Y�����P�����������uj�0�XlxVHYEB     400     1a0��7MSi�V��w~U)M݀���݇|�WN��{����'o��x1�o�l�l���^�K*�,?�^U���h�.J>Ug�Z�������\!��n�����pG3\lr� �,2�M�޶^�:KM�A�yf�F���4�ӧ�r����Pa�9�ЮbTtuѸ-��/y��nh��L;����ăO�IsN�=�,�T����0=��|����=�d�Y^S_ݜ
��Y�7�Y��x\�l�C�펗�7����IA:O�=]�J�Ie\v|R�ʳ�KOn��wJ���͌�"D;Ih���r�����h�����1읳�B|���I��v�il��3�N]3�rF��JW�:�Z�1�w�K���V�z�����i"�6�JAs�P �^,r I�2�/�>yKW��N��Dc�����K)���XlxVHYEB     400     190 ���g��}���r1;����FV�ا�\�G��7�Ğ��B�E��v�k7G�:�%���X����'�<�ѹp�]��}Y��;��Ԣ���&P9�n���r�E�$q��x�`��<�,���ܕ�>󡉑6i�l��݈��PD˾�3��&    %��d)պ5k���:��h�)5�o
���O��B�r�J,9�вG����UVMD i�B    �}ս���1u�It�    Z-Ӗ������Y>?�h?��`؞B@*oqT�Ꜣ��_�{A�<x�2_�%%X����8$`����̕推�_�b*�[i��aC�w    j�)�=��,�:s+�G���2z�ù�~½���<E���>��z/��%@�j�/�Ӻ.�W��m�k���b����,�6�XlxVHYEB     400     140}h�/
ժl�ʮ4�Ϸtz�%��L<�F�r8hL��v��Xi_�%���R�|�T������\^����6��+z������/�{����Q<���T��+<���YP�q\&���Π����Ϗ=ך�fUk?�0�¦����{:�Qn���k=�_���k\,F`�rt/P�TD1@_�I�k�f�S�H�����~Jm�����ߝ}���
��L����0x]s#]w��K²Vŀ��7Ą X�z4�3�q�_(HF"�����ƞXS�?�X�|(%ьWI�|���N�3�aB�0�5˭П=�M8qYD��xZ�L'޶XlxVHYEB     400     140/y�F��?�͉F
w��PӮ��ܧO[��O(5�^��7#��6Q}�D�v����)������U�ɡQ�����y%z��,�ZA�duz��ͳ�;_���)�ꗆ�> �<���y���)\Y}�U8�%~l��0�c�h��y��j:c趛{��f�]�s�[π@%n�}I�e�?>�i($�B�˫��    '8J6ZC��!V8���kX_?������H�-���۠���N�3���V�V��m�w\yv�ށC�Es�q�����J�����K��0��A�!L6�����<f�:�D��fcO���줥Pb�i�    �t��5EXlxVHYEB     400     150�x���9�*\�c�����K�=᫩��P�����}�4;z@��*%�U��}���b��@�$�ӕ��.ec&o��Ƙ="��L�u3>&�b��}y�tm��.��}Q���9��Đ[��:C�i�۹|ٸ�fA�������\b�0�Ì}��;d|M����lo���[`%�D�oh��3��[��g�,'`��W/y�������GM*
S�f�N]敔b�D�uE�D�=� ����+�x�_��w<�    FA�������J<z��aP���<�B�    ]`"���ج��_��~���}WT4$    U8]����Y8_��g�mə��A�4�X�ֈ�XlxVHYEB     400     140�Ru�|�ذ/0���z��X�Y
q�=2�����-�������o�\��$=훩���-��F��Rq^-�TP��M�&W�k&�     ^�w>"k�jq�v%�ؐ���&�l����J��� �X���x���M�nb[>�){�9�Sq\�������&�^J4ܮ�h E.L�/��m2�z���I�Y:'=��������R`����=��|�����xvv��@RB�4�r�=�z��R�R��:��d�u�Î��%ՁJ)MO����p;��W����m�v���+����O�K��e� {�&�Y-��O��{�N����٘yXlxVHYEB     400     1a0xe���B'�=Oǲ�P�A�/N�u�k[���4= W��0ĢS^�����6o$̽FB?��~��    1��'�-��wu�9M�|JNN���i���P��b>�ܼ�";,��v�x�!�z�S�T�͗��Ϝ]ifOv
����Zػ��4��C����~|�J�e=l�#����˿���M��<t��r2���x4��O}��aS��nI�_��}�$h��Ou�E�㟿`Hդt���'���1E�=&�LY@+�,�hbjٯfJɚ>"蔢j ���PD # �x���Lu��쓘���?�x�S���$��T�O��A��1ТrVz\��/�B��~ńf�`��������?���}��f��@5׊ާ:�,�<V�|�}]����T�&�=o�������rg�ү˘���/\�pJv^�XlxVHYEB     400     1805X# �����GoW܄c�e&2���
�bު�[�%����jT�;3U:/2���e���c!�y�Q�e2|Z��"����!�ً�ʹ�,&�),x��l���(��a�#��%ځ�HN�4m��!�~6�SZ�ʬw�~RQ��芃95�Q�^i{K�
�d
��Jݚ���T���E�����2�u�    �-��mL��>��z��wȠ ��W��3�;Yg<x����8Lܣ��t�[F�6D%��1w�'v��U����3�C��E��&}e_�ّE�mWv0`yJ�u؅� ��f�W�X�,����1hU`�����h� ���C4.�f���=���0���8f4�7ʤ��cx�s�M }����B�ݹ���Q�7�XlxVHYEB     400     140��A.��=�^/��Cn��Uivqb&�L�Ռ�.���~�̙��)�%�
�+8�ǧ,Xk��Y+hX�̢�*�|B>J�57�(�F4��c�Yuxu�d}�>G�t�g���a�m}V�4yx�"� ��B��@�E��;S������ƴ�(Cڎʐ�����6�H�/�@R�^ʒ�2��Bٖ>m<+�=vla�7�ݡ�P�ܮx��v-b����@��#ܾ�:L���U�͠-���zq�ĕo���*������)EdO&'������ym��AP(O̽��/��a*t;�)s3���~�i��sJ�X5�D��XlxVHYEB     400     170��2͖+��I���b�ҤSA���P��!uA����i�8�:}��V�`�,��@��fq���$�d{΋A�C4`c�"C���Z7|&�ੂ��s[�aPʽbe-I��*��EZ��L
�����c��G�l�%s%�ʭ�#��2g�˯:��EȳfLO���H���Y    os�����Ϫ����|;}�x'��Q|�k�����h�ƭ��Z`�CU���#V㶅X�Jl�C����0FY���Wqߗ:�,�}���˅x�
6�8l�R��\����k���\��s��<Y��YM�~�@�Y;6�b�    ��4;�xpi��D��f���n�h$�9ch���"^x0kڔNj�2�tj�E{XlxVHYEB     400     160C� 4�,z��K���    ���V�)�!�}e������G}�� ' r�c^����'L`< ��i�$XA�TҢ�$��� �k�����ňVq�<�<�58�߱_
�G��FE{����� ��@<�"'�Ry}��U�@�_e���k1�[ƈ�0���މ={����ͿD�����I����'}�P�̦�>��m)��cs���    ;���+Dr��Ǫz���HtZ˭�0);1��q|���仠�o-[��ٞ�"��(��ڳ���!�u�$3�o{cn�f@=�u[�S
D��2�����\%$��~b,)��8��p#r���ȵ�DN=0M�/�*��nXlxVHYEB     400     1a0F��#���[��-��}��J9]���y�=��$��}��-������8Z�w�����Ϩ�Qfn���"�+Y3��<�]�:��ϊ'U�2� ��n�<m��:'��ң�H�ਹ��n�& �{9������I�ꨇS�    �G}�P��4kV�Mxr��00+#\2�%b�*�.��8�+�g)�(D��d���Q~�䃟 𺀱=�)K�á���~��{h�qxJ�F7\�� )/,.�Eu�;'�@
7=@f;���}�\����N�
����-�zG��2!�����n���O46t��Ĥ��"@�������эcL8��!�@ǥ�.�xxl&���FO�������0�}��W�@��)Uґ��w�q��Y��s�_PwV��BwXlxVHYEB     400     130b�F @�X��ɮf�7���Wg�0���/�=�HV$�M���_+{������_�JR�Z�B�s�����O�O��Ϛ����JM�E���� �b��%��,�� :3ib�ԸDR�;�"2�5��~4+HDY��XɼC�mcX@�0`�=f+x'�Ոyӊg)C����b����0�s���0�HX8q�k��#�ƣ��R&���)��:â}�����l�F���luF�L���N���7�Y8;g;���p���"��,���v��;��W�㋨�P�槶��{d���rl9�?|.žXlxVHYEB     400     1a0�*�tC+���M��R�n�;�������G�4����#��f��._�f�7|�;�sd
\��ù@ʜc�z#��m�,�@0Z�����n>;��E�tl0!�.0�P�~y���ϫ(�Í� ��9+���K�%�����$�����1�s��t�:8s|�;i��������8 ���\��>�U��͎J�/�n1�4e��s��d�aŻ��mЋ=e�-��l�VŸ�/������]�3�����A�p��[�<�
N\:�������4�I'�GH���C˝|�+�����Cb}��iB-�l���m^��"7�D��rNك[���Z$<eh\�t����Ä�A��Ӓ��/    W��\w*����L�`�5�t�濟r�C"���r�?8Vc�$���    Hl�-�V00
Җ�;0�ٰ�FpXlxVHYEB     400     160�N,d�_��d�֐T��W�7�\����[[�zJ�<༆�̣�_�C����Z$�9z�#�O�]>��L1�{M&�Z��H��![s�=��X�$����땹ۅ���Hz�n�&}    >`�|H��@��{7Ւ��'����!���g ��ݓZY��s��4�^y=_h��VN�����CAnG����a�"v�{j��Ǉ��ޠ$�?ؑ^BK�+� >f��6a�#~�^J%�� &U����E�!���u�\�B�AC�Xp%���ܽH?v����ܞy��"e-�jBvi�X�-���y��2k�&�c-��v�V~oz�_.$�Y͌'s���+�+����)EY5�N$�}��CXlxVHYEB     400     150�^I�=ݑc���uS5J���uRJi�:
� �H��<���rB�db�ʘ6#�D����0��Yo��44�Z��M�E^ْ�k,��k���W|����M�`Q������iL��I��%܏iIX���    9Mcڨ�Cbɒ>W����N�(FG�L ~e,T'~F�@9��q`a% �TZd>���=ṵ��R;m��겏1��k���pZ��cj@�Ö�HAܢ��ڣ\���dق_�g1_j�����V 
�I-�h�]��k9���{���}��H��4Yw+�-�Him�$��_}:.����YEV,d�����ݶ��¹��Eo�Y�+3$%�PXlxVHYEB     400     150Ͳ�h�XZ\#��<�S�-�](�L�1�F/�p�OxG�8#��f��["A~���G��X�{�gܞŹ�[�u�n����o�ԀؼE�0�"(��N�9PX^M����M���@�����9���~������`%�-��*���c�^��A�ܷ�9ٹ��~�����Mw�j��O놥ّ���۠�tv^��Xo�KrZ�=D ֈ��4�����9P�k��@����d]��L@�d;���0w0Oa��m��cs/j��l����zp���^��Ox��?-��O?d <U�rӦ�Fh���+�L�Ad���sw0o��=�|^K�;C:<x�XlxVHYEB     400     1204t�x{�Z��9kG���j�'w�/2}���    K
�nh��8�=Ԕ�5��.ȠU5�((�Z&�c�6r �!P[�i�k�ŭ�|:j(R�){|AJT�k�##��:NLc���K$�*Q0BX^�w��v��c|q��4k�R
{�Z�H�o����x���OB�цk�B}��x*�O)|?�ܻ/�8~��9�ט���f��S_��Og����H�v���jV��ǉ�F3�澳M5E�kLa�Vt��H4���A�/֊�<��@
`9�^G��[�XlxVHYEB     400     1a0��]�87 e���� �2�����7�o�<��!mC��WNJ��4��t�h�*S�P�?G7^`Y    AY�wC���7_�"\L'����EJ�7#��Ra0m)�:"�|�7A ��;��h3���Kb��K�]�Iu:M�"J�������&ƥ�M��&�F���el� �_�Ζ��gA�&�A{��rj(���:g��Sk�:�4���x��R+�[��F���5Ѱ(��|{�bz-�n��d��θ_(��[Z����3��T/����5}l_�Q�-�s��>��㏰�J+e�ܙ�ӛ�^9�6���߰���S&l�3�� �����Y��Q*7 �̑c�h-��}�Hq���,�Vf�QW���x'֑)�1z�?U�n_�6�_���#�*߾��.D@bXlxVHYEB     400     1a0Q�W7_gtk0K�/B!�������j�è�    ���<K�;��SiIM�-o���GE�I�]P9&i�*w�\�PzK���b>����e2�~�te���|�E^U��}�4��P��~�q�ֵ=*2>�x��S�v�E����ݾ���Gn��R������<�z ���[�V��c����8�Z���{^z!����C0�s����u��������΢B�%6�s�{�.�&���?O��r�e/k�.���{�Q��l�+bsM��;r%{E��(�2�3�q�N�B�?� ����S��
yfu�@lx�\,��iQT]�ֻ�4����>`��fDq��?��[��v��dt�o���U��hiTc�
׎����n<?ǹ�:ɵBi��4����K՞h�������%ocIl�1��ؤ�<�>�zBrt�Ҷ�XlxVHYEB     400     100���S���m�m�W��;��PD��{��N�����\�gD�ބڟ�0����Jl�a̮�����r!�2�.�}��∁��%U�+��ic}+^K�}���TlԐg�F�R4�4b>�Z��ĳs�@_�%���k���    �����.}�/�T����x'�N3�d��/M���[��(�%�$A����i�fY9�/�[;RY����_iIj�Ž���8β=��g�}h�)��Ċ��|/�D���L:JӘ�óϑ�/XlxVHYEB     400      f0�%$h���)qM�x�S<jd��U�+�{�[�6r�~`��:L��4�CQ���e��9��tGտ�l1����b�v��}J��5I-8�͟�'/jyn�oWa�gZ�Ti@})�zI�8��������)=�[G�*1S�Bs&Ty�Q�;�Q_��<�'��G
��Z"
��,2�}KT�Z������1���Z��<��d���'mbm�mj�����M���*Ӥl�� ��A/ZoEp}
/����XlxVHYEB     400      f0ۚ�խi�]�d\��9F���T�2�5�Q�q󙒢    ίr�\��s��<�Ið���6�ƺ������WLPL��\��7�v'i�ĩ{dr�c�'�_�n��5t�O���'��X:y�{��}x�HHL@�d�l�^I���l&,+���lƜ/��_��.���2ߊ�/��0f�������S�6�g�ݣ�q�sǷ��w!,���(�?PO����5T�G������XlxVHYEB     400     100�+�v��K��+�!�ܨ�,�*#ժ�v�_lǲ^�[���{L��֝o9(-��s�vwFȲޕ�y��aO>5�y�k4)��!�Lq� * ��<L=���Rde}w�� �'�5�P�_.iľZng�_�g �]��k�tE�����坘C:�I����V/}��='��.��x���`c���7w!2jO&룉I��pB��]9�    h����2;��A���,�GM���k��~Z���XlxVHYEB     400      a0���78��X������۹O� �y�m�ѰA=�ƛhձfQ�g��*W#���א���c�{�E:Uת��r5��5,D�Pz�a���Ġ�mj-��is�l湫�Zw��ϻqK��r�+\��\Y��3�=z��9��G�B�-�˪ˏ�����:�縫XlxVHYEB     400      a0������    �5�d��^\l�|�����5-���G9�(��2���}��{aR܌�4v.�����X�-    ����~�U_S��>�m#�1�|^V�:'�.)����国�2j։��|i׻��?b�V�缼��m`�bL-��:�p$-�G�Ӄ�c ���m��xXlxVHYEB     400      d0��w�#_%���# (���!���xN>w��G[/�V
h�Ӏ �+[qH�FZ�v�Zy�q*�DM��%G5E�M3��eE�y�1(z��X���2c9}$VNY�    h��W�����^�j���4Y�N��;�)��}D�����*�q�5`L�0�z��S��Z�Pȧ�_i�����9�    ��s�m�.��bh�#�'\�XlxVHYEB     400      b0�{ݺ�?V1�r���3`%i!zT����5|/�    �FA�;�~��~g�}�q(Ò|c1�j-�3��3.�PbkL#�    ćf��5��>�    ��� \��q��@Og^w�n
�XR���+}�?<�BF���`���u8�n"� t��w���3��L`#eŕ�I�F*�XlxVHYEB     400     140���u�P����|E����ʮ7�VBs4�kc�Z�'�5���_��\�V��M.�)(��#��a�ʬ,���FA��^�bu��A�(���D��UT�.��g" m2���A8+�r�SL'9A�c�4����v�-h���H�Z4�YP�0A~b���Xϼ>�PB����k\���4 s�Ԙ�A]��D��FN-�    �2������Vu-��_�+�b���2��[�΢���u�����:Z�ff���
f���M�n,����E�Ybmy;f�gH5�=_��ٽ�6X����ȗ������j��0�[$P�
)�X�!��XlxVHYEB     400     120Z�S֥�H����00�9�m��6L�Qw(��;���'j��,��� �9���A�O`��La������,I�i�XH���_�ok�n��b��0����8�#��ܨq`|�"j��F.l硘���$S��ݭ��
qGTdd�496�������#*u��*JU:����J+��YH�    b+A,j�bx�;ݦj)ZV���4�Q�>�m�f�a*E������`�����D6D�    7Qq Z�4�xe�-��ֈ2e    u�"�ph���:1�Ң�G�XlxVHYEB     400     140�S�\dJՕ{.�ǌwE(�Y;�u,�nl�`��Հ��X[�c"��N�_e�]<œ�U_�R���hv��x�����D�,~��"�U�K�����n մ��J����%�(&�2�7нJ�Mͩ��4������$ғ�P�MOw0�U_�W��Ju�~P�3�����>ܾ}�! :��~�]��G�����)}0&v��A�O�;�H2��w�y�^�*���+,�c�-m�M0Yy#�,k�[US��R��fL�
��1��{Eo�B�(��qm9vb�;Lj�?�|��-�OoB����S/��mw��R猢XlxVHYEB     400     100p��c|\�VԫM��!UE��o��(���2ځնV*��m3f`��\2-������<=���E�97���]�3�@��>    ,6l�o��,�k�����x%[�7��}�<�,�����w�Tc[S��E;�0��t�T������QR�c��^�    �hv��d0�O(���Lʾ8���&�|��3g� b .��v�ʲ!�q��c��9A����5FAk�����
�����l�A̐��/    �=i��V\9`,�`7�1�XlxVHYEB     400      f0&��J��$��z��s�MWŏ&��9���
t����)&NQP��2����/[��1-�N�     ]g�4sn�!��k�4p��a�NN5B�Q�MԪc��Ð�
/������G0ֳu%��xh^m�^Q���t�����ӓ#��B�]��i(�s�$�����p��|
�@2��p��aa�V ��n�-޳*9U�/�}��Nu�´�t�w�X��,M�c���/"�}�X�s�J�p�!�fXlxVHYEB     400      e0�����|���1�h|�oZS[�fr�����Pc�B�lF�(�u[�h�_�(b�c:a��t#�{ސ�j�����P�I��5��H��    q�?o���1a��T<Ѿ�z�^��6��(��ܒbIW0���o��ȭeK��y5��'p��O�    9�QȘ�t���ߡ���|P�x2��ʋ��5Ep���C���ZTm��ƿ�<a��I"{XlxVHYEB     400      a0#S߭��<��,ڈ���|�Gm��{ɥ�����y�vV��a�2hˈ>n$H�_�At2��l�ԣ�E)G`AX1��G�l�X�ڑKmA9�!�b����j���Q�/a+�a��{Ȑ�bN�`��ĵA�l\���F�q;%�B�2(��    ��z�»�XlxVHYEB     400      a0��6*�-Y�c�ܤ����>�y���zD�0��w+��'��j)1��X���9v    ���C���c'    \;����h�ٓ��'�T�%*��=Z�n\?&:Z���i�"MMM��R�!�?;���n��S}͐ s���&s�"�5
��B�q'~�&g�:cXlxVHYEB     400      d0�i;�_�?����
��Qs�7�%�k|c�yx�u!ە�l�8�e����vU��s�}��ơ|t��݄�F��fl�z!����O������=������h����Fy)<��g9G�-�����b �=Wlb�X��a~���KP�C`��⣁r1R���/ TF?�;8/H�rs��J��V]��艾���ץ�6�G��XlxVHYEB     400      b0UIR� ����,�/�nJ�J�xϙ��'p���7� � �d�j�I��J��iZd�������*/T��ʸT�?�a/&"ē�o��I�\\���)�9v����Uμ�>�0hq/?Y?ɋ���f>n���d�~~�^~�>{ŧ��?3Q<��  �sf�#�����VIǳEx�XlxVHYEB     400     120�_g�_�a��    `QS���{�=�$���,�#��[�.�ֲmGR�'YD����D[�Q�7����`V���Dٻ�|��+��� �ײ�\�B|)��V���4�XF�D�ɮ(yӟF�4rh�/�3��LG��-�.��l�g�g���f�o�������E����'%RDJMQ +�F��͗+`���,JL���^6��&5@�_���H����<�z�'����x�    k�"Tǆ�
�">�ޛ����UMN�H�{�N�-@�H����kU;<�� _˙���P�mXlxVHYEB     400     150��3�ȱ�A{���$�4݋�!!\�0=    �T*��¾[3�]���cQ�x���#��u3Ǥ�\���y�O�J���S8��gRlp�������!�O�S��� }d,P���p>/Ro�x�{���STU<r�}N瓦�a���~[8����S"���v��{��mo��Ll�l��ю�7�6����m��a���>�6Vw��f1;҃{\mO-�-c    �RM�_9U�I���G����u�1�m_P)�p�:��o������    �m�S��95��:q-��zB5<C�b�x�O�fVB��<:�0m���|C=�5�8�W�    mx,�XlxVHYEB     400     180�$Yzj�U�*q*@�x/:�����l4B<����\��DD5|�FQ�|�*�%*�Y�H�C�J��Hg)Ⱑ��)��y�Y�j<BR;X�}��(F�����-��������n��K�evqV�X��Ʃ�9��ؿNnNi���R���B#)5ZP�����کT�����eDh��=s��پi�F    �Rh��p}&�=i�!}*2�EM��+�SI΀�e��3x��s\1s�p8����%�,jFǅ��)��
��ڮR    �_T��l�
�]��n�TN:��Iv��U���[��΁Q3����e�"��C�s*A�"��q(�

����:�    �_hs �-|�9��X[�/����$׮�f�����XlxVHYEB     400     130�$%�\-� �]4�y�W`�&Dm#�
~��    e����E&�}df/"��j�rJ+[=�s��{��D�H��1����^    ��1AM��n�ͷ#�����`�X�������i�yZ�I�=޴-��X���(��NJ��uS�wb��C��Jrp�Xl{���l�t��]�$"�H�8$O���" ����m�r��ج����8�{E�M����i�`Ӄg)�g��9���2���e1+�;�Ybv��̉B2��gm�l�����YU���շ���)����=���vِ��4�Ƙ�b�XlxVHYEB     400     170�h�����ɦ���Jg�tdac�h֬�u�� uR��|.�~��2�Z�Mw�xǥ��#�k�ȶ�=۞bK���[6Q��c�#m���e�`%e�����Xi�c���.p��s6���{'��Y�oəY���Ύ&�*b�Ae�VV����R����?�W�+';���&#�[��^
Y8�:��i�-�V��.
Ï��"�>�����R[�KРCHE�6��crax����{�D��Iclx�aN�B��5�!B�k��G T�~��q[�w��ZT���eej+�p�w���˦ҫ?b�9""����64S�+8OP�1H;�7�k�������Bk���K���7$�,���H�DDC2LT)�`��^�b���wN!XlxVHYEB     400     180(�qWm����;������ �o��F�-�"t��Z��4�p�[�G8
`A�E<��<���� ��ߔp��r�NE9��a�<\o^]^�v��f���D|Tfː�´��E�$|׋ƢJ��CU*6�ū��/7Ao��"���.�h=�U}iډ�0B����:��)]E����<ަ�H�C�NN{�@sR5�ˊ�t�q��|8#���L���j��mEP�=5���(��%��Am��e������7��n���GOz��X�����d�1#�vw��v^ ��kΞg��3��/+ci�Y6�D�    �nJ_s�Lڂ�[��.Q������<��hՑ���k�fk��0���e��*j?�΃���r� ŴȆXlxVHYEB     400     180��vk��e*�<x4T�3F���    #�����qݹs5V%qh����l �m��Ϳ�����C��^�g���b���6��E���P�X��m�{�앏P�9�{rC��!��ߔ)h�~���� �l��pM8�0�Iv��z�h�mD)fǿ�X6P�
��rd@�d�HE;�r�A*^#t�J������[�? �1t��;����a�����>"���&�    ěDN�$�����0��~�#oЦ�%9��F��V٩�����U\�Q9���3M������Paq%�l?����V�4Z.9a��P��q��ϯ5�Q���͚�cU8�i�²�T8�    ¤�W�B_��������>�w�5��( �kV���T#b��ҏ�OXlxVHYEB     400     120N��׋R2�!�eyZ7�����y?�����3��ih׎�J��@�Պ��%+���V[�E><qx�E��G�a;����7*��|�M,����    N_1N�k��y���ַQ�쥂��q(e����Z����<f�Y�����Ld'�?צ��t#�^�����ON�ի�-A��b�����X�|UlS�t zOmEta����< :�����ڳ�_��N��W�B�֣Pl��)y-ZG�g���:K�d���t�q��C"֛���C=��    J(Ѕv��XlxVHYEB     400      e0��S�6�l�-�Y�˞eEV�W%Ci�Lү�0_�����L;%����_��I|+��TO�`Ȼ!]�b���T:��#pN;g�RxP�#���D�cVE��?T��+������!�f�4G%<ć[_s�v��>�h@1"R?���¹�:��]?ŪÁ�4ʇdBm5!R�9�����i�0߯���g!�>![��NT�%�'���騂����S��@�����XlxVHYEB     400      f0�(Bݖu�Ȟ, = �Wh�v�w2#6���m,I�{�j�\K���aɈ�#��[��닭ESJ�I�z"�k����|-GO����!$�T���8����^a,]�s�:���s�������k��~�S�a+G޴V/�eܪXzqqF�ibG�-��U)+|������Hpsdd%�>���\�rL7�$��    Gԉ���h�uH������2-Y�{²��I�p�?5�XlxVHYEB     3ea      d0
f��������5�c�7�>Y1�߾X@��t䘂%�}g ~^�N�x�o�6zd��4��[c��"�&ϝUV��_�y�Օ��3���u�7�B���mA�˝�,��w԰��
?���1SdR�!���W��z�����_�����(F��7�`9�^ȬЦf�Jmt��&m��5j����k��#���T�?�g�u�'�