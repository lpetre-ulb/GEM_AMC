------------------------------------------------------------------------------------------------------------------------------------------------------
-- Company: TAMU
-- Engineer: Evaldas Juska (evaldas.juska@cern.ch, evka85@gmail.com)
-- 
-- Create Date:    12:22 2016-05-10
-- Module Name:    trigger
-- Description:    This module handles everything related to sbit cluster data (link synchronization, monitoring, local triggering, matching to L1A and reporting data to DAQ)  
------------------------------------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.numeric_std.all;

use work.gem_pkg.all;
use work.ttc_pkg.all;
use work.ipbus.all;
use work.registers.all;

entity oh_link_regs is
    generic(
        g_NUM_OF_OHs        : integer;
        g_NUM_GBTS_PER_OH   : integer
    );
    port(
        -- reset
        reset_i                 : in  std_logic;
        clk_i                   : in  std_logic;

        -- Link statuses
        gbt_link_status_arr_i   : in t_gbt_link_status_arr(g_NUM_OF_OHs * g_NUM_GBTS_PER_OH - 1 downto 0);
        vfat3_link_status_arr_i : in t_oh_vfat_link_status_arr(g_NUM_OF_OHs - 1 downto 0);

        -- Control
        vfat_mask_arr_o         : out t_std24_array(g_NUM_OF_OHs - 1 downto 0);

        -- IPbus
        ipb_reset_i             : in  std_logic;
        ipb_clk_i               : in  std_logic;
        ipb_miso_o              : out ipb_rbus;
        ipb_mosi_i              : in  ipb_wbus
    );
end oh_link_regs;

architecture oh_link_regs_arch of oh_link_regs is
    
    signal vfat_mask_arr        : t_std24_array(g_NUM_OF_OHs - 1 downto 0);
    
    ------ Register signals begin (this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py -- do not edit)
    signal regs_read_arr        : t_std32_array(REG_OH_LINKS_NUM_REGS - 1 downto 0);
    signal regs_write_arr       : t_std32_array(REG_OH_LINKS_NUM_REGS - 1 downto 0);
    signal regs_addresses       : t_std32_array(REG_OH_LINKS_NUM_REGS - 1 downto 0);
    signal regs_defaults        : t_std32_array(REG_OH_LINKS_NUM_REGS - 1 downto 0) := (others => (others => '0'));
    signal regs_read_pulse_arr  : std_logic_vector(REG_OH_LINKS_NUM_REGS - 1 downto 0);
    signal regs_write_pulse_arr : std_logic_vector(REG_OH_LINKS_NUM_REGS - 1 downto 0);
    signal regs_read_ready_arr  : std_logic_vector(REG_OH_LINKS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_write_done_arr  : std_logic_vector(REG_OH_LINKS_NUM_REGS - 1 downto 0) := (others => '1');
    signal regs_writable_arr    : std_logic_vector(REG_OH_LINKS_NUM_REGS - 1 downto 0) := (others => '0');
    ------ Register signals end ----------------------------------------------
    
begin
    
    vfat_mask_arr_o <= vfat_mask_arr;
    
    --===============================================================================================
    -- this section is generated by <gem_amc_repo_root>/scripts/generate_registers.py (do not edit) 
    --==== Registers begin ==========================================================================

    -- IPbus slave instanciation
    ipbus_slave_inst : entity work.ipbus_slave
        generic map(
           g_NUM_REGS             => REG_OH_LINKS_NUM_REGS,
           g_ADDR_HIGH_BIT        => REG_OH_LINKS_ADDRESS_MSB,
           g_ADDR_LOW_BIT         => REG_OH_LINKS_ADDRESS_LSB,
           g_USE_INDIVIDUAL_ADDRS => true
       )
       port map(
           ipb_reset_i            => ipb_reset_i,
           ipb_clk_i              => ipb_clk_i,
           ipb_mosi_i             => ipb_mosi_i,
           ipb_miso_o             => ipb_miso_o,
           usr_clk_i              => clk_i,
           regs_read_arr_i        => regs_read_arr,
           regs_write_arr_o       => regs_write_arr,
           read_pulse_arr_o       => regs_read_pulse_arr,
           write_pulse_arr_o      => regs_write_pulse_arr,
           regs_read_ready_arr_i  => regs_read_ready_arr,
           regs_write_done_arr_i  => regs_write_done_arr,
           individual_addrs_arr_i => regs_addresses,
           regs_defaults_arr_i    => regs_defaults,
           writable_regs_i        => regs_writable_arr
      );

    -- Addresses
    regs_addresses(0)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"100";
    regs_addresses(1)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"101";
    regs_addresses(2)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"110";
    regs_addresses(3)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"112";
    regs_addresses(4)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"114";
    regs_addresses(5)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"116";
    regs_addresses(6)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"118";
    regs_addresses(7)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"11a";
    regs_addresses(8)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"11c";
    regs_addresses(9)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"11e";
    regs_addresses(10)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"120";
    regs_addresses(11)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"122";
    regs_addresses(12)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"124";
    regs_addresses(13)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"126";
    regs_addresses(14)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"128";
    regs_addresses(15)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"12a";
    regs_addresses(16)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"12c";
    regs_addresses(17)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"12e";
    regs_addresses(18)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"130";
    regs_addresses(19)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"132";
    regs_addresses(20)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"134";
    regs_addresses(21)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"136";
    regs_addresses(22)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"138";
    regs_addresses(23)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"13a";
    regs_addresses(24)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"13c";
    regs_addresses(25)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"13e";
    regs_addresses(26)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"200";
    regs_addresses(27)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"201";
    regs_addresses(28)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"210";
    regs_addresses(29)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"212";
    regs_addresses(30)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"214";
    regs_addresses(31)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"216";
    regs_addresses(32)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"218";
    regs_addresses(33)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"21a";
    regs_addresses(34)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"21c";
    regs_addresses(35)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"21e";
    regs_addresses(36)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"220";
    regs_addresses(37)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"222";
    regs_addresses(38)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"224";
    regs_addresses(39)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"226";
    regs_addresses(40)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"228";
    regs_addresses(41)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"22a";
    regs_addresses(42)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"22c";
    regs_addresses(43)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"22e";
    regs_addresses(44)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"230";
    regs_addresses(45)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"232";
    regs_addresses(46)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"234";
    regs_addresses(47)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"236";
    regs_addresses(48)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"238";
    regs_addresses(49)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"23a";
    regs_addresses(50)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"23c";
    regs_addresses(51)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"23e";
    regs_addresses(52)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"300";
    regs_addresses(53)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"301";
    regs_addresses(54)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"310";
    regs_addresses(55)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"312";
    regs_addresses(56)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"314";
    regs_addresses(57)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"316";
    regs_addresses(58)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"318";
    regs_addresses(59)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"31a";
    regs_addresses(60)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"31c";
    regs_addresses(61)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"31e";
    regs_addresses(62)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"320";
    regs_addresses(63)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"322";
    regs_addresses(64)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"324";
    regs_addresses(65)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"326";
    regs_addresses(66)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"328";
    regs_addresses(67)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"32a";
    regs_addresses(68)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"32c";
    regs_addresses(69)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"32e";
    regs_addresses(70)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"330";
    regs_addresses(71)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"332";
    regs_addresses(72)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"334";
    regs_addresses(73)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"336";
    regs_addresses(74)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"338";
    regs_addresses(75)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"33a";
    regs_addresses(76)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"33c";
    regs_addresses(77)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"33e";
    regs_addresses(78)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"400";
    regs_addresses(79)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"401";
    regs_addresses(80)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"410";
    regs_addresses(81)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"412";
    regs_addresses(82)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"414";
    regs_addresses(83)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"416";
    regs_addresses(84)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"418";
    regs_addresses(85)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"41a";
    regs_addresses(86)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"41c";
    regs_addresses(87)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"41e";
    regs_addresses(88)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"420";
    regs_addresses(89)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"422";
    regs_addresses(90)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"424";
    regs_addresses(91)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"426";
    regs_addresses(92)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"428";
    regs_addresses(93)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"42a";
    regs_addresses(94)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"42c";
    regs_addresses(95)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"42e";
    regs_addresses(96)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"430";
    regs_addresses(97)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"432";
    regs_addresses(98)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"434";
    regs_addresses(99)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"436";
    regs_addresses(100)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"438";
    regs_addresses(101)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"43a";
    regs_addresses(102)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"43c";
    regs_addresses(103)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"43e";
    regs_addresses(104)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"500";
    regs_addresses(105)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"501";
    regs_addresses(106)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"510";
    regs_addresses(107)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"512";
    regs_addresses(108)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"514";
    regs_addresses(109)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"516";
    regs_addresses(110)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"518";
    regs_addresses(111)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"51a";
    regs_addresses(112)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"51c";
    regs_addresses(113)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"51e";
    regs_addresses(114)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"520";
    regs_addresses(115)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"522";
    regs_addresses(116)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"524";
    regs_addresses(117)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"526";
    regs_addresses(118)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"528";
    regs_addresses(119)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"52a";
    regs_addresses(120)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"52c";
    regs_addresses(121)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"52e";
    regs_addresses(122)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"530";
    regs_addresses(123)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"532";
    regs_addresses(124)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"534";
    regs_addresses(125)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"536";
    regs_addresses(126)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"538";
    regs_addresses(127)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"53a";
    regs_addresses(128)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"53c";
    regs_addresses(129)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"53e";
    regs_addresses(130)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"600";
    regs_addresses(131)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"601";
    regs_addresses(132)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"610";
    regs_addresses(133)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"612";
    regs_addresses(134)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"614";
    regs_addresses(135)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"616";
    regs_addresses(136)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"618";
    regs_addresses(137)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"61a";
    regs_addresses(138)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"61c";
    regs_addresses(139)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"61e";
    regs_addresses(140)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"620";
    regs_addresses(141)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"622";
    regs_addresses(142)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"624";
    regs_addresses(143)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"626";
    regs_addresses(144)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"628";
    regs_addresses(145)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"62a";
    regs_addresses(146)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"62c";
    regs_addresses(147)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"62e";
    regs_addresses(148)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"630";
    regs_addresses(149)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"632";
    regs_addresses(150)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"634";
    regs_addresses(151)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"636";
    regs_addresses(152)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"638";
    regs_addresses(153)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"63a";
    regs_addresses(154)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"63c";
    regs_addresses(155)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"63e";
    regs_addresses(156)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"700";
    regs_addresses(157)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"701";
    regs_addresses(158)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"710";
    regs_addresses(159)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"712";
    regs_addresses(160)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"714";
    regs_addresses(161)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"716";
    regs_addresses(162)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"718";
    regs_addresses(163)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"71a";
    regs_addresses(164)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"71c";
    regs_addresses(165)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"71e";
    regs_addresses(166)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"720";
    regs_addresses(167)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"722";
    regs_addresses(168)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"724";
    regs_addresses(169)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"726";
    regs_addresses(170)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"728";
    regs_addresses(171)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"72a";
    regs_addresses(172)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"72c";
    regs_addresses(173)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"72e";
    regs_addresses(174)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"730";
    regs_addresses(175)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"732";
    regs_addresses(176)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"734";
    regs_addresses(177)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"736";
    regs_addresses(178)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"738";
    regs_addresses(179)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"73a";
    regs_addresses(180)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"73c";
    regs_addresses(181)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"73e";
    regs_addresses(182)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"800";
    regs_addresses(183)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"801";
    regs_addresses(184)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"810";
    regs_addresses(185)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"812";
    regs_addresses(186)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"814";
    regs_addresses(187)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"816";
    regs_addresses(188)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"818";
    regs_addresses(189)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"81a";
    regs_addresses(190)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"81c";
    regs_addresses(191)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"81e";
    regs_addresses(192)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"820";
    regs_addresses(193)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"822";
    regs_addresses(194)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"824";
    regs_addresses(195)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"826";
    regs_addresses(196)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"828";
    regs_addresses(197)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"82a";
    regs_addresses(198)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"82c";
    regs_addresses(199)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"82e";
    regs_addresses(200)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"830";
    regs_addresses(201)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"832";
    regs_addresses(202)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"834";
    regs_addresses(203)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"836";
    regs_addresses(204)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"838";
    regs_addresses(205)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"83a";
    regs_addresses(206)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"83c";
    regs_addresses(207)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"83e";
    regs_addresses(208)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"900";
    regs_addresses(209)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"901";
    regs_addresses(210)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"910";
    regs_addresses(211)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"912";
    regs_addresses(212)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"914";
    regs_addresses(213)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"916";
    regs_addresses(214)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"918";
    regs_addresses(215)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"91a";
    regs_addresses(216)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"91c";
    regs_addresses(217)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"91e";
    regs_addresses(218)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"920";
    regs_addresses(219)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"922";
    regs_addresses(220)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"924";
    regs_addresses(221)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"926";
    regs_addresses(222)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"928";
    regs_addresses(223)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"92a";
    regs_addresses(224)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"92c";
    regs_addresses(225)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"92e";
    regs_addresses(226)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"930";
    regs_addresses(227)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"932";
    regs_addresses(228)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"934";
    regs_addresses(229)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"936";
    regs_addresses(230)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"938";
    regs_addresses(231)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"93a";
    regs_addresses(232)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"93c";
    regs_addresses(233)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"93e";
    regs_addresses(234)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a00";
    regs_addresses(235)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a01";
    regs_addresses(236)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a10";
    regs_addresses(237)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a12";
    regs_addresses(238)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a14";
    regs_addresses(239)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a16";
    regs_addresses(240)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a18";
    regs_addresses(241)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a1a";
    regs_addresses(242)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a1c";
    regs_addresses(243)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a1e";
    regs_addresses(244)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a20";
    regs_addresses(245)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a22";
    regs_addresses(246)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a24";
    regs_addresses(247)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a26";
    regs_addresses(248)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a28";
    regs_addresses(249)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a2a";
    regs_addresses(250)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a2c";
    regs_addresses(251)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a2e";
    regs_addresses(252)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a30";
    regs_addresses(253)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a32";
    regs_addresses(254)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a34";
    regs_addresses(255)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a36";
    regs_addresses(256)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a38";
    regs_addresses(257)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a3a";
    regs_addresses(258)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a3c";
    regs_addresses(259)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"a3e";
    regs_addresses(260)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b00";
    regs_addresses(261)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b01";
    regs_addresses(262)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b10";
    regs_addresses(263)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b12";
    regs_addresses(264)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b14";
    regs_addresses(265)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b16";
    regs_addresses(266)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b18";
    regs_addresses(267)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b1a";
    regs_addresses(268)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b1c";
    regs_addresses(269)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b1e";
    regs_addresses(270)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b20";
    regs_addresses(271)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b22";
    regs_addresses(272)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b24";
    regs_addresses(273)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b26";
    regs_addresses(274)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b28";
    regs_addresses(275)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b2a";
    regs_addresses(276)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b2c";
    regs_addresses(277)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b2e";
    regs_addresses(278)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b30";
    regs_addresses(279)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b32";
    regs_addresses(280)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b34";
    regs_addresses(281)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b36";
    regs_addresses(282)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b38";
    regs_addresses(283)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b3a";
    regs_addresses(284)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b3c";
    regs_addresses(285)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"b3e";
    regs_addresses(286)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c00";
    regs_addresses(287)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c01";
    regs_addresses(288)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c10";
    regs_addresses(289)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c12";
    regs_addresses(290)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c14";
    regs_addresses(291)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c16";
    regs_addresses(292)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c18";
    regs_addresses(293)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c1a";
    regs_addresses(294)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c1c";
    regs_addresses(295)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c1e";
    regs_addresses(296)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c20";
    regs_addresses(297)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c22";
    regs_addresses(298)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c24";
    regs_addresses(299)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c26";
    regs_addresses(300)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c28";
    regs_addresses(301)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c2a";
    regs_addresses(302)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c2c";
    regs_addresses(303)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c2e";
    regs_addresses(304)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c30";
    regs_addresses(305)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c32";
    regs_addresses(306)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c34";
    regs_addresses(307)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c36";
    regs_addresses(308)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c38";
    regs_addresses(309)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c3a";
    regs_addresses(310)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c3c";
    regs_addresses(311)(REG_OH_LINKS_ADDRESS_MSB downto REG_OH_LINKS_ADDRESS_LSB) <= '0' & x"c3e";

    -- Connect read signals
    regs_read_arr(0)(REG_OH_LINKS_OH0_GBT0_READY_BIT) <= gbt_link_status_arr_i(0 * g_NUM_GBTS_PER_OH + 0).gbt_rx_ready;
    regs_read_arr(0)(REG_OH_LINKS_OH0_GBT1_READY_BIT) <= gbt_link_status_arr_i(0 * g_NUM_GBTS_PER_OH + 1).gbt_rx_ready;
    regs_read_arr(0)(REG_OH_LINKS_OH0_GBT2_READY_BIT) <= gbt_link_status_arr_i(0 * g_NUM_GBTS_PER_OH + 2).gbt_rx_ready;
    regs_read_arr(0)(REG_OH_LINKS_OH0_GBT0_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(0 * g_NUM_GBTS_PER_OH + 0).gbt_rx_had_not_ready;
    regs_read_arr(0)(REG_OH_LINKS_OH0_GBT1_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(0 * g_NUM_GBTS_PER_OH + 1).gbt_rx_had_not_ready;
    regs_read_arr(0)(REG_OH_LINKS_OH0_GBT2_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(0 * g_NUM_GBTS_PER_OH + 2).gbt_rx_had_not_ready;
    regs_read_arr(0)(REG_OH_LINKS_OH0_GBT0_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(0 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_ovf;
    regs_read_arr(0)(REG_OH_LINKS_OH0_GBT1_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(0 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_ovf;
    regs_read_arr(0)(REG_OH_LINKS_OH0_GBT2_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(0 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_ovf;
    regs_read_arr(0)(REG_OH_LINKS_OH0_GBT0_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(0 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_unf;
    regs_read_arr(0)(REG_OH_LINKS_OH0_GBT1_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(0 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_unf;
    regs_read_arr(0)(REG_OH_LINKS_OH0_GBT2_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(0 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_unf;
    regs_read_arr(1)(REG_OH_LINKS_OH0_VFAT_MASK_MSB downto REG_OH_LINKS_OH0_VFAT_MASK_LSB) <= vfat_mask_arr(0);
    regs_read_arr(2)(REG_OH_LINKS_OH0_VFAT0_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(0).sync_good;
    regs_read_arr(2)(REG_OH_LINKS_OH0_VFAT0_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT0_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(0).sync_error_cnt;
    regs_read_arr(2)(REG_OH_LINKS_OH0_VFAT0_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT0_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(0).daq_event_cnt;
    regs_read_arr(2)(REG_OH_LINKS_OH0_VFAT0_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT0_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(0).daq_crc_err_cnt;
    regs_read_arr(3)(REG_OH_LINKS_OH0_VFAT1_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(1).sync_good;
    regs_read_arr(3)(REG_OH_LINKS_OH0_VFAT1_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT1_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(1).sync_error_cnt;
    regs_read_arr(3)(REG_OH_LINKS_OH0_VFAT1_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT1_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(1).daq_event_cnt;
    regs_read_arr(3)(REG_OH_LINKS_OH0_VFAT1_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT1_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(1).daq_crc_err_cnt;
    regs_read_arr(4)(REG_OH_LINKS_OH0_VFAT2_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(2).sync_good;
    regs_read_arr(4)(REG_OH_LINKS_OH0_VFAT2_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT2_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(2).sync_error_cnt;
    regs_read_arr(4)(REG_OH_LINKS_OH0_VFAT2_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT2_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(2).daq_event_cnt;
    regs_read_arr(4)(REG_OH_LINKS_OH0_VFAT2_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT2_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(2).daq_crc_err_cnt;
    regs_read_arr(5)(REG_OH_LINKS_OH0_VFAT3_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(3).sync_good;
    regs_read_arr(5)(REG_OH_LINKS_OH0_VFAT3_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT3_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(3).sync_error_cnt;
    regs_read_arr(5)(REG_OH_LINKS_OH0_VFAT3_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT3_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(3).daq_event_cnt;
    regs_read_arr(5)(REG_OH_LINKS_OH0_VFAT3_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT3_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(3).daq_crc_err_cnt;
    regs_read_arr(6)(REG_OH_LINKS_OH0_VFAT4_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(4).sync_good;
    regs_read_arr(6)(REG_OH_LINKS_OH0_VFAT4_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT4_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(4).sync_error_cnt;
    regs_read_arr(6)(REG_OH_LINKS_OH0_VFAT4_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT4_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(4).daq_event_cnt;
    regs_read_arr(6)(REG_OH_LINKS_OH0_VFAT4_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT4_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(4).daq_crc_err_cnt;
    regs_read_arr(7)(REG_OH_LINKS_OH0_VFAT5_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(5).sync_good;
    regs_read_arr(7)(REG_OH_LINKS_OH0_VFAT5_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT5_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(5).sync_error_cnt;
    regs_read_arr(7)(REG_OH_LINKS_OH0_VFAT5_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT5_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(5).daq_event_cnt;
    regs_read_arr(7)(REG_OH_LINKS_OH0_VFAT5_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT5_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(5).daq_crc_err_cnt;
    regs_read_arr(8)(REG_OH_LINKS_OH0_VFAT6_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(6).sync_good;
    regs_read_arr(8)(REG_OH_LINKS_OH0_VFAT6_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT6_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(6).sync_error_cnt;
    regs_read_arr(8)(REG_OH_LINKS_OH0_VFAT6_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT6_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(6).daq_event_cnt;
    regs_read_arr(8)(REG_OH_LINKS_OH0_VFAT6_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT6_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(6).daq_crc_err_cnt;
    regs_read_arr(9)(REG_OH_LINKS_OH0_VFAT7_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(7).sync_good;
    regs_read_arr(9)(REG_OH_LINKS_OH0_VFAT7_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT7_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(7).sync_error_cnt;
    regs_read_arr(9)(REG_OH_LINKS_OH0_VFAT7_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT7_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(7).daq_event_cnt;
    regs_read_arr(9)(REG_OH_LINKS_OH0_VFAT7_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT7_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(7).daq_crc_err_cnt;
    regs_read_arr(10)(REG_OH_LINKS_OH0_VFAT8_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(8).sync_good;
    regs_read_arr(10)(REG_OH_LINKS_OH0_VFAT8_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT8_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(8).sync_error_cnt;
    regs_read_arr(10)(REG_OH_LINKS_OH0_VFAT8_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT8_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(8).daq_event_cnt;
    regs_read_arr(10)(REG_OH_LINKS_OH0_VFAT8_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT8_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(8).daq_crc_err_cnt;
    regs_read_arr(11)(REG_OH_LINKS_OH0_VFAT9_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(9).sync_good;
    regs_read_arr(11)(REG_OH_LINKS_OH0_VFAT9_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT9_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(9).sync_error_cnt;
    regs_read_arr(11)(REG_OH_LINKS_OH0_VFAT9_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT9_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(9).daq_event_cnt;
    regs_read_arr(11)(REG_OH_LINKS_OH0_VFAT9_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT9_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(9).daq_crc_err_cnt;
    regs_read_arr(12)(REG_OH_LINKS_OH0_VFAT10_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(10).sync_good;
    regs_read_arr(12)(REG_OH_LINKS_OH0_VFAT10_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT10_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(10).sync_error_cnt;
    regs_read_arr(12)(REG_OH_LINKS_OH0_VFAT10_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT10_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(10).daq_event_cnt;
    regs_read_arr(12)(REG_OH_LINKS_OH0_VFAT10_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT10_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(10).daq_crc_err_cnt;
    regs_read_arr(13)(REG_OH_LINKS_OH0_VFAT11_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(11).sync_good;
    regs_read_arr(13)(REG_OH_LINKS_OH0_VFAT11_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT11_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(11).sync_error_cnt;
    regs_read_arr(13)(REG_OH_LINKS_OH0_VFAT11_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT11_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(11).daq_event_cnt;
    regs_read_arr(13)(REG_OH_LINKS_OH0_VFAT11_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT11_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(11).daq_crc_err_cnt;
    regs_read_arr(14)(REG_OH_LINKS_OH0_VFAT12_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(12).sync_good;
    regs_read_arr(14)(REG_OH_LINKS_OH0_VFAT12_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT12_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(12).sync_error_cnt;
    regs_read_arr(14)(REG_OH_LINKS_OH0_VFAT12_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT12_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(12).daq_event_cnt;
    regs_read_arr(14)(REG_OH_LINKS_OH0_VFAT12_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT12_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(12).daq_crc_err_cnt;
    regs_read_arr(15)(REG_OH_LINKS_OH0_VFAT13_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(13).sync_good;
    regs_read_arr(15)(REG_OH_LINKS_OH0_VFAT13_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT13_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(13).sync_error_cnt;
    regs_read_arr(15)(REG_OH_LINKS_OH0_VFAT13_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT13_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(13).daq_event_cnt;
    regs_read_arr(15)(REG_OH_LINKS_OH0_VFAT13_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT13_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(13).daq_crc_err_cnt;
    regs_read_arr(16)(REG_OH_LINKS_OH0_VFAT14_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(14).sync_good;
    regs_read_arr(16)(REG_OH_LINKS_OH0_VFAT14_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT14_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(14).sync_error_cnt;
    regs_read_arr(16)(REG_OH_LINKS_OH0_VFAT14_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT14_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(14).daq_event_cnt;
    regs_read_arr(16)(REG_OH_LINKS_OH0_VFAT14_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT14_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(14).daq_crc_err_cnt;
    regs_read_arr(17)(REG_OH_LINKS_OH0_VFAT15_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(15).sync_good;
    regs_read_arr(17)(REG_OH_LINKS_OH0_VFAT15_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT15_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(15).sync_error_cnt;
    regs_read_arr(17)(REG_OH_LINKS_OH0_VFAT15_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT15_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(15).daq_event_cnt;
    regs_read_arr(17)(REG_OH_LINKS_OH0_VFAT15_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT15_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(15).daq_crc_err_cnt;
    regs_read_arr(18)(REG_OH_LINKS_OH0_VFAT16_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(16).sync_good;
    regs_read_arr(18)(REG_OH_LINKS_OH0_VFAT16_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT16_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(16).sync_error_cnt;
    regs_read_arr(18)(REG_OH_LINKS_OH0_VFAT16_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT16_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(16).daq_event_cnt;
    regs_read_arr(18)(REG_OH_LINKS_OH0_VFAT16_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT16_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(16).daq_crc_err_cnt;
    regs_read_arr(19)(REG_OH_LINKS_OH0_VFAT17_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(17).sync_good;
    regs_read_arr(19)(REG_OH_LINKS_OH0_VFAT17_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT17_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(17).sync_error_cnt;
    regs_read_arr(19)(REG_OH_LINKS_OH0_VFAT17_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT17_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(17).daq_event_cnt;
    regs_read_arr(19)(REG_OH_LINKS_OH0_VFAT17_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT17_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(17).daq_crc_err_cnt;
    regs_read_arr(20)(REG_OH_LINKS_OH0_VFAT18_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(18).sync_good;
    regs_read_arr(20)(REG_OH_LINKS_OH0_VFAT18_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT18_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(18).sync_error_cnt;
    regs_read_arr(20)(REG_OH_LINKS_OH0_VFAT18_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT18_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(18).daq_event_cnt;
    regs_read_arr(20)(REG_OH_LINKS_OH0_VFAT18_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT18_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(18).daq_crc_err_cnt;
    regs_read_arr(21)(REG_OH_LINKS_OH0_VFAT19_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(19).sync_good;
    regs_read_arr(21)(REG_OH_LINKS_OH0_VFAT19_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT19_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(19).sync_error_cnt;
    regs_read_arr(21)(REG_OH_LINKS_OH0_VFAT19_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT19_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(19).daq_event_cnt;
    regs_read_arr(21)(REG_OH_LINKS_OH0_VFAT19_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT19_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(19).daq_crc_err_cnt;
    regs_read_arr(22)(REG_OH_LINKS_OH0_VFAT20_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(20).sync_good;
    regs_read_arr(22)(REG_OH_LINKS_OH0_VFAT20_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT20_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(20).sync_error_cnt;
    regs_read_arr(22)(REG_OH_LINKS_OH0_VFAT20_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT20_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(20).daq_event_cnt;
    regs_read_arr(22)(REG_OH_LINKS_OH0_VFAT20_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT20_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(20).daq_crc_err_cnt;
    regs_read_arr(23)(REG_OH_LINKS_OH0_VFAT21_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(21).sync_good;
    regs_read_arr(23)(REG_OH_LINKS_OH0_VFAT21_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT21_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(21).sync_error_cnt;
    regs_read_arr(23)(REG_OH_LINKS_OH0_VFAT21_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT21_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(21).daq_event_cnt;
    regs_read_arr(23)(REG_OH_LINKS_OH0_VFAT21_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT21_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(21).daq_crc_err_cnt;
    regs_read_arr(24)(REG_OH_LINKS_OH0_VFAT22_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(22).sync_good;
    regs_read_arr(24)(REG_OH_LINKS_OH0_VFAT22_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT22_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(22).sync_error_cnt;
    regs_read_arr(24)(REG_OH_LINKS_OH0_VFAT22_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT22_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(22).daq_event_cnt;
    regs_read_arr(24)(REG_OH_LINKS_OH0_VFAT22_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT22_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(22).daq_crc_err_cnt;
    regs_read_arr(25)(REG_OH_LINKS_OH0_VFAT23_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(0)(23).sync_good;
    regs_read_arr(25)(REG_OH_LINKS_OH0_VFAT23_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT23_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(0)(23).sync_error_cnt;
    regs_read_arr(25)(REG_OH_LINKS_OH0_VFAT23_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH0_VFAT23_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(0)(23).daq_event_cnt;
    regs_read_arr(25)(REG_OH_LINKS_OH0_VFAT23_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH0_VFAT23_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(0)(23).daq_crc_err_cnt;
    regs_read_arr(26)(REG_OH_LINKS_OH1_GBT0_READY_BIT) <= gbt_link_status_arr_i(1 * g_NUM_GBTS_PER_OH + 0).gbt_rx_ready;
    regs_read_arr(26)(REG_OH_LINKS_OH1_GBT1_READY_BIT) <= gbt_link_status_arr_i(1 * g_NUM_GBTS_PER_OH + 1).gbt_rx_ready;
    regs_read_arr(26)(REG_OH_LINKS_OH1_GBT2_READY_BIT) <= gbt_link_status_arr_i(1 * g_NUM_GBTS_PER_OH + 2).gbt_rx_ready;
    regs_read_arr(26)(REG_OH_LINKS_OH1_GBT0_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(1 * g_NUM_GBTS_PER_OH + 0).gbt_rx_had_not_ready;
    regs_read_arr(26)(REG_OH_LINKS_OH1_GBT1_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(1 * g_NUM_GBTS_PER_OH + 1).gbt_rx_had_not_ready;
    regs_read_arr(26)(REG_OH_LINKS_OH1_GBT2_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(1 * g_NUM_GBTS_PER_OH + 2).gbt_rx_had_not_ready;
    regs_read_arr(26)(REG_OH_LINKS_OH1_GBT0_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(1 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_ovf;
    regs_read_arr(26)(REG_OH_LINKS_OH1_GBT1_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(1 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_ovf;
    regs_read_arr(26)(REG_OH_LINKS_OH1_GBT2_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(1 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_ovf;
    regs_read_arr(26)(REG_OH_LINKS_OH1_GBT0_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(1 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_unf;
    regs_read_arr(26)(REG_OH_LINKS_OH1_GBT1_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(1 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_unf;
    regs_read_arr(26)(REG_OH_LINKS_OH1_GBT2_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(1 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_unf;
    regs_read_arr(27)(REG_OH_LINKS_OH1_VFAT_MASK_MSB downto REG_OH_LINKS_OH1_VFAT_MASK_LSB) <= vfat_mask_arr(1);
    regs_read_arr(28)(REG_OH_LINKS_OH1_VFAT0_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(0).sync_good;
    regs_read_arr(28)(REG_OH_LINKS_OH1_VFAT0_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT0_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(0).sync_error_cnt;
    regs_read_arr(28)(REG_OH_LINKS_OH1_VFAT0_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT0_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(0).daq_event_cnt;
    regs_read_arr(28)(REG_OH_LINKS_OH1_VFAT0_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT0_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(0).daq_crc_err_cnt;
    regs_read_arr(29)(REG_OH_LINKS_OH1_VFAT1_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(1).sync_good;
    regs_read_arr(29)(REG_OH_LINKS_OH1_VFAT1_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT1_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(1).sync_error_cnt;
    regs_read_arr(29)(REG_OH_LINKS_OH1_VFAT1_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT1_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(1).daq_event_cnt;
    regs_read_arr(29)(REG_OH_LINKS_OH1_VFAT1_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT1_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(1).daq_crc_err_cnt;
    regs_read_arr(30)(REG_OH_LINKS_OH1_VFAT2_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(2).sync_good;
    regs_read_arr(30)(REG_OH_LINKS_OH1_VFAT2_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT2_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(2).sync_error_cnt;
    regs_read_arr(30)(REG_OH_LINKS_OH1_VFAT2_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT2_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(2).daq_event_cnt;
    regs_read_arr(30)(REG_OH_LINKS_OH1_VFAT2_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT2_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(2).daq_crc_err_cnt;
    regs_read_arr(31)(REG_OH_LINKS_OH1_VFAT3_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(3).sync_good;
    regs_read_arr(31)(REG_OH_LINKS_OH1_VFAT3_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT3_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(3).sync_error_cnt;
    regs_read_arr(31)(REG_OH_LINKS_OH1_VFAT3_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT3_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(3).daq_event_cnt;
    regs_read_arr(31)(REG_OH_LINKS_OH1_VFAT3_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT3_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(3).daq_crc_err_cnt;
    regs_read_arr(32)(REG_OH_LINKS_OH1_VFAT4_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(4).sync_good;
    regs_read_arr(32)(REG_OH_LINKS_OH1_VFAT4_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT4_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(4).sync_error_cnt;
    regs_read_arr(32)(REG_OH_LINKS_OH1_VFAT4_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT4_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(4).daq_event_cnt;
    regs_read_arr(32)(REG_OH_LINKS_OH1_VFAT4_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT4_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(4).daq_crc_err_cnt;
    regs_read_arr(33)(REG_OH_LINKS_OH1_VFAT5_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(5).sync_good;
    regs_read_arr(33)(REG_OH_LINKS_OH1_VFAT5_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT5_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(5).sync_error_cnt;
    regs_read_arr(33)(REG_OH_LINKS_OH1_VFAT5_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT5_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(5).daq_event_cnt;
    regs_read_arr(33)(REG_OH_LINKS_OH1_VFAT5_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT5_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(5).daq_crc_err_cnt;
    regs_read_arr(34)(REG_OH_LINKS_OH1_VFAT6_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(6).sync_good;
    regs_read_arr(34)(REG_OH_LINKS_OH1_VFAT6_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT6_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(6).sync_error_cnt;
    regs_read_arr(34)(REG_OH_LINKS_OH1_VFAT6_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT6_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(6).daq_event_cnt;
    regs_read_arr(34)(REG_OH_LINKS_OH1_VFAT6_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT6_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(6).daq_crc_err_cnt;
    regs_read_arr(35)(REG_OH_LINKS_OH1_VFAT7_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(7).sync_good;
    regs_read_arr(35)(REG_OH_LINKS_OH1_VFAT7_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT7_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(7).sync_error_cnt;
    regs_read_arr(35)(REG_OH_LINKS_OH1_VFAT7_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT7_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(7).daq_event_cnt;
    regs_read_arr(35)(REG_OH_LINKS_OH1_VFAT7_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT7_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(7).daq_crc_err_cnt;
    regs_read_arr(36)(REG_OH_LINKS_OH1_VFAT8_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(8).sync_good;
    regs_read_arr(36)(REG_OH_LINKS_OH1_VFAT8_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT8_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(8).sync_error_cnt;
    regs_read_arr(36)(REG_OH_LINKS_OH1_VFAT8_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT8_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(8).daq_event_cnt;
    regs_read_arr(36)(REG_OH_LINKS_OH1_VFAT8_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT8_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(8).daq_crc_err_cnt;
    regs_read_arr(37)(REG_OH_LINKS_OH1_VFAT9_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(9).sync_good;
    regs_read_arr(37)(REG_OH_LINKS_OH1_VFAT9_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT9_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(9).sync_error_cnt;
    regs_read_arr(37)(REG_OH_LINKS_OH1_VFAT9_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT9_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(9).daq_event_cnt;
    regs_read_arr(37)(REG_OH_LINKS_OH1_VFAT9_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT9_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(9).daq_crc_err_cnt;
    regs_read_arr(38)(REG_OH_LINKS_OH1_VFAT10_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(10).sync_good;
    regs_read_arr(38)(REG_OH_LINKS_OH1_VFAT10_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT10_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(10).sync_error_cnt;
    regs_read_arr(38)(REG_OH_LINKS_OH1_VFAT10_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT10_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(10).daq_event_cnt;
    regs_read_arr(38)(REG_OH_LINKS_OH1_VFAT10_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT10_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(10).daq_crc_err_cnt;
    regs_read_arr(39)(REG_OH_LINKS_OH1_VFAT11_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(11).sync_good;
    regs_read_arr(39)(REG_OH_LINKS_OH1_VFAT11_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT11_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(11).sync_error_cnt;
    regs_read_arr(39)(REG_OH_LINKS_OH1_VFAT11_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT11_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(11).daq_event_cnt;
    regs_read_arr(39)(REG_OH_LINKS_OH1_VFAT11_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT11_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(11).daq_crc_err_cnt;
    regs_read_arr(40)(REG_OH_LINKS_OH1_VFAT12_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(12).sync_good;
    regs_read_arr(40)(REG_OH_LINKS_OH1_VFAT12_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT12_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(12).sync_error_cnt;
    regs_read_arr(40)(REG_OH_LINKS_OH1_VFAT12_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT12_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(12).daq_event_cnt;
    regs_read_arr(40)(REG_OH_LINKS_OH1_VFAT12_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT12_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(12).daq_crc_err_cnt;
    regs_read_arr(41)(REG_OH_LINKS_OH1_VFAT13_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(13).sync_good;
    regs_read_arr(41)(REG_OH_LINKS_OH1_VFAT13_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT13_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(13).sync_error_cnt;
    regs_read_arr(41)(REG_OH_LINKS_OH1_VFAT13_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT13_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(13).daq_event_cnt;
    regs_read_arr(41)(REG_OH_LINKS_OH1_VFAT13_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT13_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(13).daq_crc_err_cnt;
    regs_read_arr(42)(REG_OH_LINKS_OH1_VFAT14_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(14).sync_good;
    regs_read_arr(42)(REG_OH_LINKS_OH1_VFAT14_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT14_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(14).sync_error_cnt;
    regs_read_arr(42)(REG_OH_LINKS_OH1_VFAT14_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT14_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(14).daq_event_cnt;
    regs_read_arr(42)(REG_OH_LINKS_OH1_VFAT14_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT14_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(14).daq_crc_err_cnt;
    regs_read_arr(43)(REG_OH_LINKS_OH1_VFAT15_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(15).sync_good;
    regs_read_arr(43)(REG_OH_LINKS_OH1_VFAT15_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT15_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(15).sync_error_cnt;
    regs_read_arr(43)(REG_OH_LINKS_OH1_VFAT15_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT15_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(15).daq_event_cnt;
    regs_read_arr(43)(REG_OH_LINKS_OH1_VFAT15_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT15_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(15).daq_crc_err_cnt;
    regs_read_arr(44)(REG_OH_LINKS_OH1_VFAT16_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(16).sync_good;
    regs_read_arr(44)(REG_OH_LINKS_OH1_VFAT16_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT16_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(16).sync_error_cnt;
    regs_read_arr(44)(REG_OH_LINKS_OH1_VFAT16_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT16_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(16).daq_event_cnt;
    regs_read_arr(44)(REG_OH_LINKS_OH1_VFAT16_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT16_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(16).daq_crc_err_cnt;
    regs_read_arr(45)(REG_OH_LINKS_OH1_VFAT17_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(17).sync_good;
    regs_read_arr(45)(REG_OH_LINKS_OH1_VFAT17_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT17_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(17).sync_error_cnt;
    regs_read_arr(45)(REG_OH_LINKS_OH1_VFAT17_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT17_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(17).daq_event_cnt;
    regs_read_arr(45)(REG_OH_LINKS_OH1_VFAT17_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT17_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(17).daq_crc_err_cnt;
    regs_read_arr(46)(REG_OH_LINKS_OH1_VFAT18_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(18).sync_good;
    regs_read_arr(46)(REG_OH_LINKS_OH1_VFAT18_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT18_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(18).sync_error_cnt;
    regs_read_arr(46)(REG_OH_LINKS_OH1_VFAT18_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT18_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(18).daq_event_cnt;
    regs_read_arr(46)(REG_OH_LINKS_OH1_VFAT18_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT18_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(18).daq_crc_err_cnt;
    regs_read_arr(47)(REG_OH_LINKS_OH1_VFAT19_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(19).sync_good;
    regs_read_arr(47)(REG_OH_LINKS_OH1_VFAT19_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT19_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(19).sync_error_cnt;
    regs_read_arr(47)(REG_OH_LINKS_OH1_VFAT19_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT19_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(19).daq_event_cnt;
    regs_read_arr(47)(REG_OH_LINKS_OH1_VFAT19_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT19_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(19).daq_crc_err_cnt;
    regs_read_arr(48)(REG_OH_LINKS_OH1_VFAT20_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(20).sync_good;
    regs_read_arr(48)(REG_OH_LINKS_OH1_VFAT20_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT20_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(20).sync_error_cnt;
    regs_read_arr(48)(REG_OH_LINKS_OH1_VFAT20_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT20_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(20).daq_event_cnt;
    regs_read_arr(48)(REG_OH_LINKS_OH1_VFAT20_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT20_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(20).daq_crc_err_cnt;
    regs_read_arr(49)(REG_OH_LINKS_OH1_VFAT21_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(21).sync_good;
    regs_read_arr(49)(REG_OH_LINKS_OH1_VFAT21_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT21_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(21).sync_error_cnt;
    regs_read_arr(49)(REG_OH_LINKS_OH1_VFAT21_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT21_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(21).daq_event_cnt;
    regs_read_arr(49)(REG_OH_LINKS_OH1_VFAT21_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT21_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(21).daq_crc_err_cnt;
    regs_read_arr(50)(REG_OH_LINKS_OH1_VFAT22_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(22).sync_good;
    regs_read_arr(50)(REG_OH_LINKS_OH1_VFAT22_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT22_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(22).sync_error_cnt;
    regs_read_arr(50)(REG_OH_LINKS_OH1_VFAT22_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT22_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(22).daq_event_cnt;
    regs_read_arr(50)(REG_OH_LINKS_OH1_VFAT22_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT22_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(22).daq_crc_err_cnt;
    regs_read_arr(51)(REG_OH_LINKS_OH1_VFAT23_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(1)(23).sync_good;
    regs_read_arr(51)(REG_OH_LINKS_OH1_VFAT23_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT23_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(1)(23).sync_error_cnt;
    regs_read_arr(51)(REG_OH_LINKS_OH1_VFAT23_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH1_VFAT23_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(1)(23).daq_event_cnt;
    regs_read_arr(51)(REG_OH_LINKS_OH1_VFAT23_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH1_VFAT23_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(1)(23).daq_crc_err_cnt;
    regs_read_arr(52)(REG_OH_LINKS_OH2_GBT0_READY_BIT) <= gbt_link_status_arr_i(2 * g_NUM_GBTS_PER_OH + 0).gbt_rx_ready;
    regs_read_arr(52)(REG_OH_LINKS_OH2_GBT1_READY_BIT) <= gbt_link_status_arr_i(2 * g_NUM_GBTS_PER_OH + 1).gbt_rx_ready;
    regs_read_arr(52)(REG_OH_LINKS_OH2_GBT2_READY_BIT) <= gbt_link_status_arr_i(2 * g_NUM_GBTS_PER_OH + 2).gbt_rx_ready;
    regs_read_arr(52)(REG_OH_LINKS_OH2_GBT0_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(2 * g_NUM_GBTS_PER_OH + 0).gbt_rx_had_not_ready;
    regs_read_arr(52)(REG_OH_LINKS_OH2_GBT1_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(2 * g_NUM_GBTS_PER_OH + 1).gbt_rx_had_not_ready;
    regs_read_arr(52)(REG_OH_LINKS_OH2_GBT2_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(2 * g_NUM_GBTS_PER_OH + 2).gbt_rx_had_not_ready;
    regs_read_arr(52)(REG_OH_LINKS_OH2_GBT0_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(2 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_ovf;
    regs_read_arr(52)(REG_OH_LINKS_OH2_GBT1_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(2 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_ovf;
    regs_read_arr(52)(REG_OH_LINKS_OH2_GBT2_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(2 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_ovf;
    regs_read_arr(52)(REG_OH_LINKS_OH2_GBT0_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(2 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_unf;
    regs_read_arr(52)(REG_OH_LINKS_OH2_GBT1_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(2 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_unf;
    regs_read_arr(52)(REG_OH_LINKS_OH2_GBT2_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(2 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_unf;
    regs_read_arr(53)(REG_OH_LINKS_OH2_VFAT_MASK_MSB downto REG_OH_LINKS_OH2_VFAT_MASK_LSB) <= vfat_mask_arr(2);
    regs_read_arr(54)(REG_OH_LINKS_OH2_VFAT0_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(0).sync_good;
    regs_read_arr(54)(REG_OH_LINKS_OH2_VFAT0_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT0_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(0).sync_error_cnt;
    regs_read_arr(54)(REG_OH_LINKS_OH2_VFAT0_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT0_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(0).daq_event_cnt;
    regs_read_arr(54)(REG_OH_LINKS_OH2_VFAT0_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT0_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(0).daq_crc_err_cnt;
    regs_read_arr(55)(REG_OH_LINKS_OH2_VFAT1_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(1).sync_good;
    regs_read_arr(55)(REG_OH_LINKS_OH2_VFAT1_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT1_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(1).sync_error_cnt;
    regs_read_arr(55)(REG_OH_LINKS_OH2_VFAT1_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT1_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(1).daq_event_cnt;
    regs_read_arr(55)(REG_OH_LINKS_OH2_VFAT1_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT1_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(1).daq_crc_err_cnt;
    regs_read_arr(56)(REG_OH_LINKS_OH2_VFAT2_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(2).sync_good;
    regs_read_arr(56)(REG_OH_LINKS_OH2_VFAT2_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT2_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(2).sync_error_cnt;
    regs_read_arr(56)(REG_OH_LINKS_OH2_VFAT2_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT2_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(2).daq_event_cnt;
    regs_read_arr(56)(REG_OH_LINKS_OH2_VFAT2_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT2_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(2).daq_crc_err_cnt;
    regs_read_arr(57)(REG_OH_LINKS_OH2_VFAT3_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(3).sync_good;
    regs_read_arr(57)(REG_OH_LINKS_OH2_VFAT3_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT3_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(3).sync_error_cnt;
    regs_read_arr(57)(REG_OH_LINKS_OH2_VFAT3_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT3_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(3).daq_event_cnt;
    regs_read_arr(57)(REG_OH_LINKS_OH2_VFAT3_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT3_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(3).daq_crc_err_cnt;
    regs_read_arr(58)(REG_OH_LINKS_OH2_VFAT4_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(4).sync_good;
    regs_read_arr(58)(REG_OH_LINKS_OH2_VFAT4_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT4_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(4).sync_error_cnt;
    regs_read_arr(58)(REG_OH_LINKS_OH2_VFAT4_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT4_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(4).daq_event_cnt;
    regs_read_arr(58)(REG_OH_LINKS_OH2_VFAT4_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT4_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(4).daq_crc_err_cnt;
    regs_read_arr(59)(REG_OH_LINKS_OH2_VFAT5_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(5).sync_good;
    regs_read_arr(59)(REG_OH_LINKS_OH2_VFAT5_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT5_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(5).sync_error_cnt;
    regs_read_arr(59)(REG_OH_LINKS_OH2_VFAT5_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT5_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(5).daq_event_cnt;
    regs_read_arr(59)(REG_OH_LINKS_OH2_VFAT5_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT5_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(5).daq_crc_err_cnt;
    regs_read_arr(60)(REG_OH_LINKS_OH2_VFAT6_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(6).sync_good;
    regs_read_arr(60)(REG_OH_LINKS_OH2_VFAT6_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT6_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(6).sync_error_cnt;
    regs_read_arr(60)(REG_OH_LINKS_OH2_VFAT6_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT6_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(6).daq_event_cnt;
    regs_read_arr(60)(REG_OH_LINKS_OH2_VFAT6_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT6_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(6).daq_crc_err_cnt;
    regs_read_arr(61)(REG_OH_LINKS_OH2_VFAT7_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(7).sync_good;
    regs_read_arr(61)(REG_OH_LINKS_OH2_VFAT7_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT7_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(7).sync_error_cnt;
    regs_read_arr(61)(REG_OH_LINKS_OH2_VFAT7_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT7_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(7).daq_event_cnt;
    regs_read_arr(61)(REG_OH_LINKS_OH2_VFAT7_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT7_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(7).daq_crc_err_cnt;
    regs_read_arr(62)(REG_OH_LINKS_OH2_VFAT8_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(8).sync_good;
    regs_read_arr(62)(REG_OH_LINKS_OH2_VFAT8_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT8_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(8).sync_error_cnt;
    regs_read_arr(62)(REG_OH_LINKS_OH2_VFAT8_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT8_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(8).daq_event_cnt;
    regs_read_arr(62)(REG_OH_LINKS_OH2_VFAT8_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT8_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(8).daq_crc_err_cnt;
    regs_read_arr(63)(REG_OH_LINKS_OH2_VFAT9_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(9).sync_good;
    regs_read_arr(63)(REG_OH_LINKS_OH2_VFAT9_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT9_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(9).sync_error_cnt;
    regs_read_arr(63)(REG_OH_LINKS_OH2_VFAT9_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT9_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(9).daq_event_cnt;
    regs_read_arr(63)(REG_OH_LINKS_OH2_VFAT9_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT9_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(9).daq_crc_err_cnt;
    regs_read_arr(64)(REG_OH_LINKS_OH2_VFAT10_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(10).sync_good;
    regs_read_arr(64)(REG_OH_LINKS_OH2_VFAT10_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT10_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(10).sync_error_cnt;
    regs_read_arr(64)(REG_OH_LINKS_OH2_VFAT10_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT10_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(10).daq_event_cnt;
    regs_read_arr(64)(REG_OH_LINKS_OH2_VFAT10_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT10_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(10).daq_crc_err_cnt;
    regs_read_arr(65)(REG_OH_LINKS_OH2_VFAT11_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(11).sync_good;
    regs_read_arr(65)(REG_OH_LINKS_OH2_VFAT11_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT11_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(11).sync_error_cnt;
    regs_read_arr(65)(REG_OH_LINKS_OH2_VFAT11_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT11_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(11).daq_event_cnt;
    regs_read_arr(65)(REG_OH_LINKS_OH2_VFAT11_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT11_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(11).daq_crc_err_cnt;
    regs_read_arr(66)(REG_OH_LINKS_OH2_VFAT12_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(12).sync_good;
    regs_read_arr(66)(REG_OH_LINKS_OH2_VFAT12_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT12_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(12).sync_error_cnt;
    regs_read_arr(66)(REG_OH_LINKS_OH2_VFAT12_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT12_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(12).daq_event_cnt;
    regs_read_arr(66)(REG_OH_LINKS_OH2_VFAT12_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT12_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(12).daq_crc_err_cnt;
    regs_read_arr(67)(REG_OH_LINKS_OH2_VFAT13_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(13).sync_good;
    regs_read_arr(67)(REG_OH_LINKS_OH2_VFAT13_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT13_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(13).sync_error_cnt;
    regs_read_arr(67)(REG_OH_LINKS_OH2_VFAT13_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT13_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(13).daq_event_cnt;
    regs_read_arr(67)(REG_OH_LINKS_OH2_VFAT13_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT13_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(13).daq_crc_err_cnt;
    regs_read_arr(68)(REG_OH_LINKS_OH2_VFAT14_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(14).sync_good;
    regs_read_arr(68)(REG_OH_LINKS_OH2_VFAT14_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT14_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(14).sync_error_cnt;
    regs_read_arr(68)(REG_OH_LINKS_OH2_VFAT14_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT14_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(14).daq_event_cnt;
    regs_read_arr(68)(REG_OH_LINKS_OH2_VFAT14_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT14_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(14).daq_crc_err_cnt;
    regs_read_arr(69)(REG_OH_LINKS_OH2_VFAT15_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(15).sync_good;
    regs_read_arr(69)(REG_OH_LINKS_OH2_VFAT15_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT15_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(15).sync_error_cnt;
    regs_read_arr(69)(REG_OH_LINKS_OH2_VFAT15_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT15_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(15).daq_event_cnt;
    regs_read_arr(69)(REG_OH_LINKS_OH2_VFAT15_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT15_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(15).daq_crc_err_cnt;
    regs_read_arr(70)(REG_OH_LINKS_OH2_VFAT16_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(16).sync_good;
    regs_read_arr(70)(REG_OH_LINKS_OH2_VFAT16_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT16_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(16).sync_error_cnt;
    regs_read_arr(70)(REG_OH_LINKS_OH2_VFAT16_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT16_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(16).daq_event_cnt;
    regs_read_arr(70)(REG_OH_LINKS_OH2_VFAT16_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT16_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(16).daq_crc_err_cnt;
    regs_read_arr(71)(REG_OH_LINKS_OH2_VFAT17_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(17).sync_good;
    regs_read_arr(71)(REG_OH_LINKS_OH2_VFAT17_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT17_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(17).sync_error_cnt;
    regs_read_arr(71)(REG_OH_LINKS_OH2_VFAT17_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT17_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(17).daq_event_cnt;
    regs_read_arr(71)(REG_OH_LINKS_OH2_VFAT17_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT17_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(17).daq_crc_err_cnt;
    regs_read_arr(72)(REG_OH_LINKS_OH2_VFAT18_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(18).sync_good;
    regs_read_arr(72)(REG_OH_LINKS_OH2_VFAT18_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT18_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(18).sync_error_cnt;
    regs_read_arr(72)(REG_OH_LINKS_OH2_VFAT18_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT18_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(18).daq_event_cnt;
    regs_read_arr(72)(REG_OH_LINKS_OH2_VFAT18_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT18_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(18).daq_crc_err_cnt;
    regs_read_arr(73)(REG_OH_LINKS_OH2_VFAT19_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(19).sync_good;
    regs_read_arr(73)(REG_OH_LINKS_OH2_VFAT19_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT19_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(19).sync_error_cnt;
    regs_read_arr(73)(REG_OH_LINKS_OH2_VFAT19_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT19_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(19).daq_event_cnt;
    regs_read_arr(73)(REG_OH_LINKS_OH2_VFAT19_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT19_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(19).daq_crc_err_cnt;
    regs_read_arr(74)(REG_OH_LINKS_OH2_VFAT20_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(20).sync_good;
    regs_read_arr(74)(REG_OH_LINKS_OH2_VFAT20_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT20_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(20).sync_error_cnt;
    regs_read_arr(74)(REG_OH_LINKS_OH2_VFAT20_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT20_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(20).daq_event_cnt;
    regs_read_arr(74)(REG_OH_LINKS_OH2_VFAT20_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT20_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(20).daq_crc_err_cnt;
    regs_read_arr(75)(REG_OH_LINKS_OH2_VFAT21_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(21).sync_good;
    regs_read_arr(75)(REG_OH_LINKS_OH2_VFAT21_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT21_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(21).sync_error_cnt;
    regs_read_arr(75)(REG_OH_LINKS_OH2_VFAT21_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT21_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(21).daq_event_cnt;
    regs_read_arr(75)(REG_OH_LINKS_OH2_VFAT21_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT21_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(21).daq_crc_err_cnt;
    regs_read_arr(76)(REG_OH_LINKS_OH2_VFAT22_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(22).sync_good;
    regs_read_arr(76)(REG_OH_LINKS_OH2_VFAT22_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT22_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(22).sync_error_cnt;
    regs_read_arr(76)(REG_OH_LINKS_OH2_VFAT22_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT22_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(22).daq_event_cnt;
    regs_read_arr(76)(REG_OH_LINKS_OH2_VFAT22_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT22_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(22).daq_crc_err_cnt;
    regs_read_arr(77)(REG_OH_LINKS_OH2_VFAT23_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(2)(23).sync_good;
    regs_read_arr(77)(REG_OH_LINKS_OH2_VFAT23_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT23_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(2)(23).sync_error_cnt;
    regs_read_arr(77)(REG_OH_LINKS_OH2_VFAT23_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH2_VFAT23_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(2)(23).daq_event_cnt;
    regs_read_arr(77)(REG_OH_LINKS_OH2_VFAT23_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH2_VFAT23_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(2)(23).daq_crc_err_cnt;
    regs_read_arr(78)(REG_OH_LINKS_OH3_GBT0_READY_BIT) <= gbt_link_status_arr_i(3 * g_NUM_GBTS_PER_OH + 0).gbt_rx_ready;
    regs_read_arr(78)(REG_OH_LINKS_OH3_GBT1_READY_BIT) <= gbt_link_status_arr_i(3 * g_NUM_GBTS_PER_OH + 1).gbt_rx_ready;
    regs_read_arr(78)(REG_OH_LINKS_OH3_GBT2_READY_BIT) <= gbt_link_status_arr_i(3 * g_NUM_GBTS_PER_OH + 2).gbt_rx_ready;
    regs_read_arr(78)(REG_OH_LINKS_OH3_GBT0_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(3 * g_NUM_GBTS_PER_OH + 0).gbt_rx_had_not_ready;
    regs_read_arr(78)(REG_OH_LINKS_OH3_GBT1_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(3 * g_NUM_GBTS_PER_OH + 1).gbt_rx_had_not_ready;
    regs_read_arr(78)(REG_OH_LINKS_OH3_GBT2_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(3 * g_NUM_GBTS_PER_OH + 2).gbt_rx_had_not_ready;
    regs_read_arr(78)(REG_OH_LINKS_OH3_GBT0_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(3 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_ovf;
    regs_read_arr(78)(REG_OH_LINKS_OH3_GBT1_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(3 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_ovf;
    regs_read_arr(78)(REG_OH_LINKS_OH3_GBT2_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(3 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_ovf;
    regs_read_arr(78)(REG_OH_LINKS_OH3_GBT0_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(3 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_unf;
    regs_read_arr(78)(REG_OH_LINKS_OH3_GBT1_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(3 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_unf;
    regs_read_arr(78)(REG_OH_LINKS_OH3_GBT2_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(3 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_unf;
    regs_read_arr(79)(REG_OH_LINKS_OH3_VFAT_MASK_MSB downto REG_OH_LINKS_OH3_VFAT_MASK_LSB) <= vfat_mask_arr(3);
    regs_read_arr(80)(REG_OH_LINKS_OH3_VFAT0_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(0).sync_good;
    regs_read_arr(80)(REG_OH_LINKS_OH3_VFAT0_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT0_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(0).sync_error_cnt;
    regs_read_arr(80)(REG_OH_LINKS_OH3_VFAT0_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT0_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(0).daq_event_cnt;
    regs_read_arr(80)(REG_OH_LINKS_OH3_VFAT0_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT0_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(0).daq_crc_err_cnt;
    regs_read_arr(81)(REG_OH_LINKS_OH3_VFAT1_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(1).sync_good;
    regs_read_arr(81)(REG_OH_LINKS_OH3_VFAT1_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT1_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(1).sync_error_cnt;
    regs_read_arr(81)(REG_OH_LINKS_OH3_VFAT1_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT1_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(1).daq_event_cnt;
    regs_read_arr(81)(REG_OH_LINKS_OH3_VFAT1_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT1_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(1).daq_crc_err_cnt;
    regs_read_arr(82)(REG_OH_LINKS_OH3_VFAT2_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(2).sync_good;
    regs_read_arr(82)(REG_OH_LINKS_OH3_VFAT2_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT2_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(2).sync_error_cnt;
    regs_read_arr(82)(REG_OH_LINKS_OH3_VFAT2_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT2_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(2).daq_event_cnt;
    regs_read_arr(82)(REG_OH_LINKS_OH3_VFAT2_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT2_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(2).daq_crc_err_cnt;
    regs_read_arr(83)(REG_OH_LINKS_OH3_VFAT3_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(3).sync_good;
    regs_read_arr(83)(REG_OH_LINKS_OH3_VFAT3_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT3_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(3).sync_error_cnt;
    regs_read_arr(83)(REG_OH_LINKS_OH3_VFAT3_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT3_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(3).daq_event_cnt;
    regs_read_arr(83)(REG_OH_LINKS_OH3_VFAT3_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT3_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(3).daq_crc_err_cnt;
    regs_read_arr(84)(REG_OH_LINKS_OH3_VFAT4_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(4).sync_good;
    regs_read_arr(84)(REG_OH_LINKS_OH3_VFAT4_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT4_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(4).sync_error_cnt;
    regs_read_arr(84)(REG_OH_LINKS_OH3_VFAT4_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT4_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(4).daq_event_cnt;
    regs_read_arr(84)(REG_OH_LINKS_OH3_VFAT4_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT4_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(4).daq_crc_err_cnt;
    regs_read_arr(85)(REG_OH_LINKS_OH3_VFAT5_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(5).sync_good;
    regs_read_arr(85)(REG_OH_LINKS_OH3_VFAT5_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT5_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(5).sync_error_cnt;
    regs_read_arr(85)(REG_OH_LINKS_OH3_VFAT5_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT5_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(5).daq_event_cnt;
    regs_read_arr(85)(REG_OH_LINKS_OH3_VFAT5_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT5_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(5).daq_crc_err_cnt;
    regs_read_arr(86)(REG_OH_LINKS_OH3_VFAT6_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(6).sync_good;
    regs_read_arr(86)(REG_OH_LINKS_OH3_VFAT6_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT6_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(6).sync_error_cnt;
    regs_read_arr(86)(REG_OH_LINKS_OH3_VFAT6_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT6_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(6).daq_event_cnt;
    regs_read_arr(86)(REG_OH_LINKS_OH3_VFAT6_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT6_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(6).daq_crc_err_cnt;
    regs_read_arr(87)(REG_OH_LINKS_OH3_VFAT7_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(7).sync_good;
    regs_read_arr(87)(REG_OH_LINKS_OH3_VFAT7_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT7_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(7).sync_error_cnt;
    regs_read_arr(87)(REG_OH_LINKS_OH3_VFAT7_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT7_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(7).daq_event_cnt;
    regs_read_arr(87)(REG_OH_LINKS_OH3_VFAT7_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT7_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(7).daq_crc_err_cnt;
    regs_read_arr(88)(REG_OH_LINKS_OH3_VFAT8_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(8).sync_good;
    regs_read_arr(88)(REG_OH_LINKS_OH3_VFAT8_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT8_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(8).sync_error_cnt;
    regs_read_arr(88)(REG_OH_LINKS_OH3_VFAT8_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT8_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(8).daq_event_cnt;
    regs_read_arr(88)(REG_OH_LINKS_OH3_VFAT8_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT8_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(8).daq_crc_err_cnt;
    regs_read_arr(89)(REG_OH_LINKS_OH3_VFAT9_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(9).sync_good;
    regs_read_arr(89)(REG_OH_LINKS_OH3_VFAT9_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT9_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(9).sync_error_cnt;
    regs_read_arr(89)(REG_OH_LINKS_OH3_VFAT9_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT9_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(9).daq_event_cnt;
    regs_read_arr(89)(REG_OH_LINKS_OH3_VFAT9_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT9_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(9).daq_crc_err_cnt;
    regs_read_arr(90)(REG_OH_LINKS_OH3_VFAT10_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(10).sync_good;
    regs_read_arr(90)(REG_OH_LINKS_OH3_VFAT10_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT10_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(10).sync_error_cnt;
    regs_read_arr(90)(REG_OH_LINKS_OH3_VFAT10_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT10_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(10).daq_event_cnt;
    regs_read_arr(90)(REG_OH_LINKS_OH3_VFAT10_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT10_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(10).daq_crc_err_cnt;
    regs_read_arr(91)(REG_OH_LINKS_OH3_VFAT11_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(11).sync_good;
    regs_read_arr(91)(REG_OH_LINKS_OH3_VFAT11_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT11_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(11).sync_error_cnt;
    regs_read_arr(91)(REG_OH_LINKS_OH3_VFAT11_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT11_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(11).daq_event_cnt;
    regs_read_arr(91)(REG_OH_LINKS_OH3_VFAT11_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT11_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(11).daq_crc_err_cnt;
    regs_read_arr(92)(REG_OH_LINKS_OH3_VFAT12_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(12).sync_good;
    regs_read_arr(92)(REG_OH_LINKS_OH3_VFAT12_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT12_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(12).sync_error_cnt;
    regs_read_arr(92)(REG_OH_LINKS_OH3_VFAT12_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT12_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(12).daq_event_cnt;
    regs_read_arr(92)(REG_OH_LINKS_OH3_VFAT12_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT12_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(12).daq_crc_err_cnt;
    regs_read_arr(93)(REG_OH_LINKS_OH3_VFAT13_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(13).sync_good;
    regs_read_arr(93)(REG_OH_LINKS_OH3_VFAT13_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT13_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(13).sync_error_cnt;
    regs_read_arr(93)(REG_OH_LINKS_OH3_VFAT13_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT13_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(13).daq_event_cnt;
    regs_read_arr(93)(REG_OH_LINKS_OH3_VFAT13_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT13_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(13).daq_crc_err_cnt;
    regs_read_arr(94)(REG_OH_LINKS_OH3_VFAT14_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(14).sync_good;
    regs_read_arr(94)(REG_OH_LINKS_OH3_VFAT14_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT14_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(14).sync_error_cnt;
    regs_read_arr(94)(REG_OH_LINKS_OH3_VFAT14_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT14_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(14).daq_event_cnt;
    regs_read_arr(94)(REG_OH_LINKS_OH3_VFAT14_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT14_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(14).daq_crc_err_cnt;
    regs_read_arr(95)(REG_OH_LINKS_OH3_VFAT15_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(15).sync_good;
    regs_read_arr(95)(REG_OH_LINKS_OH3_VFAT15_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT15_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(15).sync_error_cnt;
    regs_read_arr(95)(REG_OH_LINKS_OH3_VFAT15_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT15_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(15).daq_event_cnt;
    regs_read_arr(95)(REG_OH_LINKS_OH3_VFAT15_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT15_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(15).daq_crc_err_cnt;
    regs_read_arr(96)(REG_OH_LINKS_OH3_VFAT16_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(16).sync_good;
    regs_read_arr(96)(REG_OH_LINKS_OH3_VFAT16_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT16_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(16).sync_error_cnt;
    regs_read_arr(96)(REG_OH_LINKS_OH3_VFAT16_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT16_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(16).daq_event_cnt;
    regs_read_arr(96)(REG_OH_LINKS_OH3_VFAT16_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT16_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(16).daq_crc_err_cnt;
    regs_read_arr(97)(REG_OH_LINKS_OH3_VFAT17_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(17).sync_good;
    regs_read_arr(97)(REG_OH_LINKS_OH3_VFAT17_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT17_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(17).sync_error_cnt;
    regs_read_arr(97)(REG_OH_LINKS_OH3_VFAT17_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT17_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(17).daq_event_cnt;
    regs_read_arr(97)(REG_OH_LINKS_OH3_VFAT17_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT17_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(17).daq_crc_err_cnt;
    regs_read_arr(98)(REG_OH_LINKS_OH3_VFAT18_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(18).sync_good;
    regs_read_arr(98)(REG_OH_LINKS_OH3_VFAT18_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT18_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(18).sync_error_cnt;
    regs_read_arr(98)(REG_OH_LINKS_OH3_VFAT18_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT18_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(18).daq_event_cnt;
    regs_read_arr(98)(REG_OH_LINKS_OH3_VFAT18_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT18_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(18).daq_crc_err_cnt;
    regs_read_arr(99)(REG_OH_LINKS_OH3_VFAT19_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(19).sync_good;
    regs_read_arr(99)(REG_OH_LINKS_OH3_VFAT19_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT19_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(19).sync_error_cnt;
    regs_read_arr(99)(REG_OH_LINKS_OH3_VFAT19_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT19_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(19).daq_event_cnt;
    regs_read_arr(99)(REG_OH_LINKS_OH3_VFAT19_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT19_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(19).daq_crc_err_cnt;
    regs_read_arr(100)(REG_OH_LINKS_OH3_VFAT20_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(20).sync_good;
    regs_read_arr(100)(REG_OH_LINKS_OH3_VFAT20_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT20_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(20).sync_error_cnt;
    regs_read_arr(100)(REG_OH_LINKS_OH3_VFAT20_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT20_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(20).daq_event_cnt;
    regs_read_arr(100)(REG_OH_LINKS_OH3_VFAT20_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT20_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(20).daq_crc_err_cnt;
    regs_read_arr(101)(REG_OH_LINKS_OH3_VFAT21_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(21).sync_good;
    regs_read_arr(101)(REG_OH_LINKS_OH3_VFAT21_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT21_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(21).sync_error_cnt;
    regs_read_arr(101)(REG_OH_LINKS_OH3_VFAT21_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT21_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(21).daq_event_cnt;
    regs_read_arr(101)(REG_OH_LINKS_OH3_VFAT21_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT21_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(21).daq_crc_err_cnt;
    regs_read_arr(102)(REG_OH_LINKS_OH3_VFAT22_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(22).sync_good;
    regs_read_arr(102)(REG_OH_LINKS_OH3_VFAT22_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT22_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(22).sync_error_cnt;
    regs_read_arr(102)(REG_OH_LINKS_OH3_VFAT22_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT22_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(22).daq_event_cnt;
    regs_read_arr(102)(REG_OH_LINKS_OH3_VFAT22_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT22_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(22).daq_crc_err_cnt;
    regs_read_arr(103)(REG_OH_LINKS_OH3_VFAT23_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(3)(23).sync_good;
    regs_read_arr(103)(REG_OH_LINKS_OH3_VFAT23_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT23_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(3)(23).sync_error_cnt;
    regs_read_arr(103)(REG_OH_LINKS_OH3_VFAT23_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH3_VFAT23_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(3)(23).daq_event_cnt;
    regs_read_arr(103)(REG_OH_LINKS_OH3_VFAT23_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH3_VFAT23_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(3)(23).daq_crc_err_cnt;
    regs_read_arr(104)(REG_OH_LINKS_OH4_GBT0_READY_BIT) <= gbt_link_status_arr_i(4 * g_NUM_GBTS_PER_OH + 0).gbt_rx_ready;
    regs_read_arr(104)(REG_OH_LINKS_OH4_GBT1_READY_BIT) <= gbt_link_status_arr_i(4 * g_NUM_GBTS_PER_OH + 1).gbt_rx_ready;
    regs_read_arr(104)(REG_OH_LINKS_OH4_GBT2_READY_BIT) <= gbt_link_status_arr_i(4 * g_NUM_GBTS_PER_OH + 2).gbt_rx_ready;
    regs_read_arr(104)(REG_OH_LINKS_OH4_GBT0_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(4 * g_NUM_GBTS_PER_OH + 0).gbt_rx_had_not_ready;
    regs_read_arr(104)(REG_OH_LINKS_OH4_GBT1_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(4 * g_NUM_GBTS_PER_OH + 1).gbt_rx_had_not_ready;
    regs_read_arr(104)(REG_OH_LINKS_OH4_GBT2_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(4 * g_NUM_GBTS_PER_OH + 2).gbt_rx_had_not_ready;
    regs_read_arr(104)(REG_OH_LINKS_OH4_GBT0_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(4 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_ovf;
    regs_read_arr(104)(REG_OH_LINKS_OH4_GBT1_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(4 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_ovf;
    regs_read_arr(104)(REG_OH_LINKS_OH4_GBT2_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(4 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_ovf;
    regs_read_arr(104)(REG_OH_LINKS_OH4_GBT0_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(4 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_unf;
    regs_read_arr(104)(REG_OH_LINKS_OH4_GBT1_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(4 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_unf;
    regs_read_arr(104)(REG_OH_LINKS_OH4_GBT2_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(4 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_unf;
    regs_read_arr(105)(REG_OH_LINKS_OH4_VFAT_MASK_MSB downto REG_OH_LINKS_OH4_VFAT_MASK_LSB) <= vfat_mask_arr(4);
    regs_read_arr(106)(REG_OH_LINKS_OH4_VFAT0_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(0).sync_good;
    regs_read_arr(106)(REG_OH_LINKS_OH4_VFAT0_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT0_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(0).sync_error_cnt;
    regs_read_arr(106)(REG_OH_LINKS_OH4_VFAT0_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT0_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(0).daq_event_cnt;
    regs_read_arr(106)(REG_OH_LINKS_OH4_VFAT0_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT0_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(0).daq_crc_err_cnt;
    regs_read_arr(107)(REG_OH_LINKS_OH4_VFAT1_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(1).sync_good;
    regs_read_arr(107)(REG_OH_LINKS_OH4_VFAT1_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT1_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(1).sync_error_cnt;
    regs_read_arr(107)(REG_OH_LINKS_OH4_VFAT1_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT1_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(1).daq_event_cnt;
    regs_read_arr(107)(REG_OH_LINKS_OH4_VFAT1_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT1_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(1).daq_crc_err_cnt;
    regs_read_arr(108)(REG_OH_LINKS_OH4_VFAT2_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(2).sync_good;
    regs_read_arr(108)(REG_OH_LINKS_OH4_VFAT2_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT2_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(2).sync_error_cnt;
    regs_read_arr(108)(REG_OH_LINKS_OH4_VFAT2_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT2_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(2).daq_event_cnt;
    regs_read_arr(108)(REG_OH_LINKS_OH4_VFAT2_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT2_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(2).daq_crc_err_cnt;
    regs_read_arr(109)(REG_OH_LINKS_OH4_VFAT3_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(3).sync_good;
    regs_read_arr(109)(REG_OH_LINKS_OH4_VFAT3_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT3_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(3).sync_error_cnt;
    regs_read_arr(109)(REG_OH_LINKS_OH4_VFAT3_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT3_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(3).daq_event_cnt;
    regs_read_arr(109)(REG_OH_LINKS_OH4_VFAT3_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT3_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(3).daq_crc_err_cnt;
    regs_read_arr(110)(REG_OH_LINKS_OH4_VFAT4_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(4).sync_good;
    regs_read_arr(110)(REG_OH_LINKS_OH4_VFAT4_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT4_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(4).sync_error_cnt;
    regs_read_arr(110)(REG_OH_LINKS_OH4_VFAT4_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT4_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(4).daq_event_cnt;
    regs_read_arr(110)(REG_OH_LINKS_OH4_VFAT4_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT4_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(4).daq_crc_err_cnt;
    regs_read_arr(111)(REG_OH_LINKS_OH4_VFAT5_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(5).sync_good;
    regs_read_arr(111)(REG_OH_LINKS_OH4_VFAT5_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT5_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(5).sync_error_cnt;
    regs_read_arr(111)(REG_OH_LINKS_OH4_VFAT5_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT5_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(5).daq_event_cnt;
    regs_read_arr(111)(REG_OH_LINKS_OH4_VFAT5_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT5_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(5).daq_crc_err_cnt;
    regs_read_arr(112)(REG_OH_LINKS_OH4_VFAT6_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(6).sync_good;
    regs_read_arr(112)(REG_OH_LINKS_OH4_VFAT6_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT6_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(6).sync_error_cnt;
    regs_read_arr(112)(REG_OH_LINKS_OH4_VFAT6_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT6_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(6).daq_event_cnt;
    regs_read_arr(112)(REG_OH_LINKS_OH4_VFAT6_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT6_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(6).daq_crc_err_cnt;
    regs_read_arr(113)(REG_OH_LINKS_OH4_VFAT7_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(7).sync_good;
    regs_read_arr(113)(REG_OH_LINKS_OH4_VFAT7_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT7_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(7).sync_error_cnt;
    regs_read_arr(113)(REG_OH_LINKS_OH4_VFAT7_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT7_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(7).daq_event_cnt;
    regs_read_arr(113)(REG_OH_LINKS_OH4_VFAT7_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT7_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(7).daq_crc_err_cnt;
    regs_read_arr(114)(REG_OH_LINKS_OH4_VFAT8_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(8).sync_good;
    regs_read_arr(114)(REG_OH_LINKS_OH4_VFAT8_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT8_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(8).sync_error_cnt;
    regs_read_arr(114)(REG_OH_LINKS_OH4_VFAT8_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT8_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(8).daq_event_cnt;
    regs_read_arr(114)(REG_OH_LINKS_OH4_VFAT8_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT8_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(8).daq_crc_err_cnt;
    regs_read_arr(115)(REG_OH_LINKS_OH4_VFAT9_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(9).sync_good;
    regs_read_arr(115)(REG_OH_LINKS_OH4_VFAT9_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT9_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(9).sync_error_cnt;
    regs_read_arr(115)(REG_OH_LINKS_OH4_VFAT9_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT9_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(9).daq_event_cnt;
    regs_read_arr(115)(REG_OH_LINKS_OH4_VFAT9_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT9_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(9).daq_crc_err_cnt;
    regs_read_arr(116)(REG_OH_LINKS_OH4_VFAT10_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(10).sync_good;
    regs_read_arr(116)(REG_OH_LINKS_OH4_VFAT10_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT10_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(10).sync_error_cnt;
    regs_read_arr(116)(REG_OH_LINKS_OH4_VFAT10_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT10_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(10).daq_event_cnt;
    regs_read_arr(116)(REG_OH_LINKS_OH4_VFAT10_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT10_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(10).daq_crc_err_cnt;
    regs_read_arr(117)(REG_OH_LINKS_OH4_VFAT11_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(11).sync_good;
    regs_read_arr(117)(REG_OH_LINKS_OH4_VFAT11_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT11_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(11).sync_error_cnt;
    regs_read_arr(117)(REG_OH_LINKS_OH4_VFAT11_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT11_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(11).daq_event_cnt;
    regs_read_arr(117)(REG_OH_LINKS_OH4_VFAT11_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT11_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(11).daq_crc_err_cnt;
    regs_read_arr(118)(REG_OH_LINKS_OH4_VFAT12_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(12).sync_good;
    regs_read_arr(118)(REG_OH_LINKS_OH4_VFAT12_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT12_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(12).sync_error_cnt;
    regs_read_arr(118)(REG_OH_LINKS_OH4_VFAT12_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT12_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(12).daq_event_cnt;
    regs_read_arr(118)(REG_OH_LINKS_OH4_VFAT12_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT12_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(12).daq_crc_err_cnt;
    regs_read_arr(119)(REG_OH_LINKS_OH4_VFAT13_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(13).sync_good;
    regs_read_arr(119)(REG_OH_LINKS_OH4_VFAT13_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT13_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(13).sync_error_cnt;
    regs_read_arr(119)(REG_OH_LINKS_OH4_VFAT13_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT13_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(13).daq_event_cnt;
    regs_read_arr(119)(REG_OH_LINKS_OH4_VFAT13_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT13_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(13).daq_crc_err_cnt;
    regs_read_arr(120)(REG_OH_LINKS_OH4_VFAT14_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(14).sync_good;
    regs_read_arr(120)(REG_OH_LINKS_OH4_VFAT14_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT14_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(14).sync_error_cnt;
    regs_read_arr(120)(REG_OH_LINKS_OH4_VFAT14_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT14_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(14).daq_event_cnt;
    regs_read_arr(120)(REG_OH_LINKS_OH4_VFAT14_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT14_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(14).daq_crc_err_cnt;
    regs_read_arr(121)(REG_OH_LINKS_OH4_VFAT15_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(15).sync_good;
    regs_read_arr(121)(REG_OH_LINKS_OH4_VFAT15_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT15_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(15).sync_error_cnt;
    regs_read_arr(121)(REG_OH_LINKS_OH4_VFAT15_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT15_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(15).daq_event_cnt;
    regs_read_arr(121)(REG_OH_LINKS_OH4_VFAT15_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT15_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(15).daq_crc_err_cnt;
    regs_read_arr(122)(REG_OH_LINKS_OH4_VFAT16_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(16).sync_good;
    regs_read_arr(122)(REG_OH_LINKS_OH4_VFAT16_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT16_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(16).sync_error_cnt;
    regs_read_arr(122)(REG_OH_LINKS_OH4_VFAT16_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT16_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(16).daq_event_cnt;
    regs_read_arr(122)(REG_OH_LINKS_OH4_VFAT16_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT16_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(16).daq_crc_err_cnt;
    regs_read_arr(123)(REG_OH_LINKS_OH4_VFAT17_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(17).sync_good;
    regs_read_arr(123)(REG_OH_LINKS_OH4_VFAT17_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT17_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(17).sync_error_cnt;
    regs_read_arr(123)(REG_OH_LINKS_OH4_VFAT17_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT17_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(17).daq_event_cnt;
    regs_read_arr(123)(REG_OH_LINKS_OH4_VFAT17_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT17_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(17).daq_crc_err_cnt;
    regs_read_arr(124)(REG_OH_LINKS_OH4_VFAT18_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(18).sync_good;
    regs_read_arr(124)(REG_OH_LINKS_OH4_VFAT18_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT18_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(18).sync_error_cnt;
    regs_read_arr(124)(REG_OH_LINKS_OH4_VFAT18_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT18_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(18).daq_event_cnt;
    regs_read_arr(124)(REG_OH_LINKS_OH4_VFAT18_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT18_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(18).daq_crc_err_cnt;
    regs_read_arr(125)(REG_OH_LINKS_OH4_VFAT19_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(19).sync_good;
    regs_read_arr(125)(REG_OH_LINKS_OH4_VFAT19_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT19_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(19).sync_error_cnt;
    regs_read_arr(125)(REG_OH_LINKS_OH4_VFAT19_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT19_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(19).daq_event_cnt;
    regs_read_arr(125)(REG_OH_LINKS_OH4_VFAT19_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT19_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(19).daq_crc_err_cnt;
    regs_read_arr(126)(REG_OH_LINKS_OH4_VFAT20_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(20).sync_good;
    regs_read_arr(126)(REG_OH_LINKS_OH4_VFAT20_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT20_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(20).sync_error_cnt;
    regs_read_arr(126)(REG_OH_LINKS_OH4_VFAT20_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT20_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(20).daq_event_cnt;
    regs_read_arr(126)(REG_OH_LINKS_OH4_VFAT20_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT20_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(20).daq_crc_err_cnt;
    regs_read_arr(127)(REG_OH_LINKS_OH4_VFAT21_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(21).sync_good;
    regs_read_arr(127)(REG_OH_LINKS_OH4_VFAT21_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT21_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(21).sync_error_cnt;
    regs_read_arr(127)(REG_OH_LINKS_OH4_VFAT21_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT21_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(21).daq_event_cnt;
    regs_read_arr(127)(REG_OH_LINKS_OH4_VFAT21_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT21_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(21).daq_crc_err_cnt;
    regs_read_arr(128)(REG_OH_LINKS_OH4_VFAT22_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(22).sync_good;
    regs_read_arr(128)(REG_OH_LINKS_OH4_VFAT22_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT22_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(22).sync_error_cnt;
    regs_read_arr(128)(REG_OH_LINKS_OH4_VFAT22_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT22_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(22).daq_event_cnt;
    regs_read_arr(128)(REG_OH_LINKS_OH4_VFAT22_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT22_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(22).daq_crc_err_cnt;
    regs_read_arr(129)(REG_OH_LINKS_OH4_VFAT23_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(4)(23).sync_good;
    regs_read_arr(129)(REG_OH_LINKS_OH4_VFAT23_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT23_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(4)(23).sync_error_cnt;
    regs_read_arr(129)(REG_OH_LINKS_OH4_VFAT23_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH4_VFAT23_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(4)(23).daq_event_cnt;
    regs_read_arr(129)(REG_OH_LINKS_OH4_VFAT23_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH4_VFAT23_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(4)(23).daq_crc_err_cnt;
    regs_read_arr(130)(REG_OH_LINKS_OH5_GBT0_READY_BIT) <= gbt_link_status_arr_i(5 * g_NUM_GBTS_PER_OH + 0).gbt_rx_ready;
    regs_read_arr(130)(REG_OH_LINKS_OH5_GBT1_READY_BIT) <= gbt_link_status_arr_i(5 * g_NUM_GBTS_PER_OH + 1).gbt_rx_ready;
    regs_read_arr(130)(REG_OH_LINKS_OH5_GBT2_READY_BIT) <= gbt_link_status_arr_i(5 * g_NUM_GBTS_PER_OH + 2).gbt_rx_ready;
    regs_read_arr(130)(REG_OH_LINKS_OH5_GBT0_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(5 * g_NUM_GBTS_PER_OH + 0).gbt_rx_had_not_ready;
    regs_read_arr(130)(REG_OH_LINKS_OH5_GBT1_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(5 * g_NUM_GBTS_PER_OH + 1).gbt_rx_had_not_ready;
    regs_read_arr(130)(REG_OH_LINKS_OH5_GBT2_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(5 * g_NUM_GBTS_PER_OH + 2).gbt_rx_had_not_ready;
    regs_read_arr(130)(REG_OH_LINKS_OH5_GBT0_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(5 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_ovf;
    regs_read_arr(130)(REG_OH_LINKS_OH5_GBT1_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(5 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_ovf;
    regs_read_arr(130)(REG_OH_LINKS_OH5_GBT2_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(5 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_ovf;
    regs_read_arr(130)(REG_OH_LINKS_OH5_GBT0_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(5 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_unf;
    regs_read_arr(130)(REG_OH_LINKS_OH5_GBT1_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(5 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_unf;
    regs_read_arr(130)(REG_OH_LINKS_OH5_GBT2_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(5 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_unf;
    regs_read_arr(131)(REG_OH_LINKS_OH5_VFAT_MASK_MSB downto REG_OH_LINKS_OH5_VFAT_MASK_LSB) <= vfat_mask_arr(5);
    regs_read_arr(132)(REG_OH_LINKS_OH5_VFAT0_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(0).sync_good;
    regs_read_arr(132)(REG_OH_LINKS_OH5_VFAT0_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT0_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(0).sync_error_cnt;
    regs_read_arr(132)(REG_OH_LINKS_OH5_VFAT0_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT0_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(0).daq_event_cnt;
    regs_read_arr(132)(REG_OH_LINKS_OH5_VFAT0_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT0_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(0).daq_crc_err_cnt;
    regs_read_arr(133)(REG_OH_LINKS_OH5_VFAT1_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(1).sync_good;
    regs_read_arr(133)(REG_OH_LINKS_OH5_VFAT1_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT1_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(1).sync_error_cnt;
    regs_read_arr(133)(REG_OH_LINKS_OH5_VFAT1_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT1_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(1).daq_event_cnt;
    regs_read_arr(133)(REG_OH_LINKS_OH5_VFAT1_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT1_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(1).daq_crc_err_cnt;
    regs_read_arr(134)(REG_OH_LINKS_OH5_VFAT2_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(2).sync_good;
    regs_read_arr(134)(REG_OH_LINKS_OH5_VFAT2_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT2_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(2).sync_error_cnt;
    regs_read_arr(134)(REG_OH_LINKS_OH5_VFAT2_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT2_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(2).daq_event_cnt;
    regs_read_arr(134)(REG_OH_LINKS_OH5_VFAT2_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT2_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(2).daq_crc_err_cnt;
    regs_read_arr(135)(REG_OH_LINKS_OH5_VFAT3_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(3).sync_good;
    regs_read_arr(135)(REG_OH_LINKS_OH5_VFAT3_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT3_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(3).sync_error_cnt;
    regs_read_arr(135)(REG_OH_LINKS_OH5_VFAT3_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT3_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(3).daq_event_cnt;
    regs_read_arr(135)(REG_OH_LINKS_OH5_VFAT3_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT3_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(3).daq_crc_err_cnt;
    regs_read_arr(136)(REG_OH_LINKS_OH5_VFAT4_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(4).sync_good;
    regs_read_arr(136)(REG_OH_LINKS_OH5_VFAT4_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT4_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(4).sync_error_cnt;
    regs_read_arr(136)(REG_OH_LINKS_OH5_VFAT4_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT4_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(4).daq_event_cnt;
    regs_read_arr(136)(REG_OH_LINKS_OH5_VFAT4_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT4_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(4).daq_crc_err_cnt;
    regs_read_arr(137)(REG_OH_LINKS_OH5_VFAT5_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(5).sync_good;
    regs_read_arr(137)(REG_OH_LINKS_OH5_VFAT5_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT5_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(5).sync_error_cnt;
    regs_read_arr(137)(REG_OH_LINKS_OH5_VFAT5_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT5_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(5).daq_event_cnt;
    regs_read_arr(137)(REG_OH_LINKS_OH5_VFAT5_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT5_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(5).daq_crc_err_cnt;
    regs_read_arr(138)(REG_OH_LINKS_OH5_VFAT6_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(6).sync_good;
    regs_read_arr(138)(REG_OH_LINKS_OH5_VFAT6_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT6_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(6).sync_error_cnt;
    regs_read_arr(138)(REG_OH_LINKS_OH5_VFAT6_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT6_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(6).daq_event_cnt;
    regs_read_arr(138)(REG_OH_LINKS_OH5_VFAT6_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT6_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(6).daq_crc_err_cnt;
    regs_read_arr(139)(REG_OH_LINKS_OH5_VFAT7_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(7).sync_good;
    regs_read_arr(139)(REG_OH_LINKS_OH5_VFAT7_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT7_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(7).sync_error_cnt;
    regs_read_arr(139)(REG_OH_LINKS_OH5_VFAT7_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT7_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(7).daq_event_cnt;
    regs_read_arr(139)(REG_OH_LINKS_OH5_VFAT7_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT7_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(7).daq_crc_err_cnt;
    regs_read_arr(140)(REG_OH_LINKS_OH5_VFAT8_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(8).sync_good;
    regs_read_arr(140)(REG_OH_LINKS_OH5_VFAT8_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT8_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(8).sync_error_cnt;
    regs_read_arr(140)(REG_OH_LINKS_OH5_VFAT8_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT8_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(8).daq_event_cnt;
    regs_read_arr(140)(REG_OH_LINKS_OH5_VFAT8_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT8_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(8).daq_crc_err_cnt;
    regs_read_arr(141)(REG_OH_LINKS_OH5_VFAT9_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(9).sync_good;
    regs_read_arr(141)(REG_OH_LINKS_OH5_VFAT9_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT9_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(9).sync_error_cnt;
    regs_read_arr(141)(REG_OH_LINKS_OH5_VFAT9_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT9_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(9).daq_event_cnt;
    regs_read_arr(141)(REG_OH_LINKS_OH5_VFAT9_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT9_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(9).daq_crc_err_cnt;
    regs_read_arr(142)(REG_OH_LINKS_OH5_VFAT10_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(10).sync_good;
    regs_read_arr(142)(REG_OH_LINKS_OH5_VFAT10_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT10_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(10).sync_error_cnt;
    regs_read_arr(142)(REG_OH_LINKS_OH5_VFAT10_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT10_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(10).daq_event_cnt;
    regs_read_arr(142)(REG_OH_LINKS_OH5_VFAT10_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT10_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(10).daq_crc_err_cnt;
    regs_read_arr(143)(REG_OH_LINKS_OH5_VFAT11_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(11).sync_good;
    regs_read_arr(143)(REG_OH_LINKS_OH5_VFAT11_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT11_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(11).sync_error_cnt;
    regs_read_arr(143)(REG_OH_LINKS_OH5_VFAT11_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT11_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(11).daq_event_cnt;
    regs_read_arr(143)(REG_OH_LINKS_OH5_VFAT11_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT11_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(11).daq_crc_err_cnt;
    regs_read_arr(144)(REG_OH_LINKS_OH5_VFAT12_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(12).sync_good;
    regs_read_arr(144)(REG_OH_LINKS_OH5_VFAT12_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT12_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(12).sync_error_cnt;
    regs_read_arr(144)(REG_OH_LINKS_OH5_VFAT12_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT12_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(12).daq_event_cnt;
    regs_read_arr(144)(REG_OH_LINKS_OH5_VFAT12_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT12_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(12).daq_crc_err_cnt;
    regs_read_arr(145)(REG_OH_LINKS_OH5_VFAT13_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(13).sync_good;
    regs_read_arr(145)(REG_OH_LINKS_OH5_VFAT13_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT13_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(13).sync_error_cnt;
    regs_read_arr(145)(REG_OH_LINKS_OH5_VFAT13_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT13_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(13).daq_event_cnt;
    regs_read_arr(145)(REG_OH_LINKS_OH5_VFAT13_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT13_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(13).daq_crc_err_cnt;
    regs_read_arr(146)(REG_OH_LINKS_OH5_VFAT14_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(14).sync_good;
    regs_read_arr(146)(REG_OH_LINKS_OH5_VFAT14_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT14_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(14).sync_error_cnt;
    regs_read_arr(146)(REG_OH_LINKS_OH5_VFAT14_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT14_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(14).daq_event_cnt;
    regs_read_arr(146)(REG_OH_LINKS_OH5_VFAT14_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT14_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(14).daq_crc_err_cnt;
    regs_read_arr(147)(REG_OH_LINKS_OH5_VFAT15_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(15).sync_good;
    regs_read_arr(147)(REG_OH_LINKS_OH5_VFAT15_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT15_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(15).sync_error_cnt;
    regs_read_arr(147)(REG_OH_LINKS_OH5_VFAT15_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT15_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(15).daq_event_cnt;
    regs_read_arr(147)(REG_OH_LINKS_OH5_VFAT15_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT15_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(15).daq_crc_err_cnt;
    regs_read_arr(148)(REG_OH_LINKS_OH5_VFAT16_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(16).sync_good;
    regs_read_arr(148)(REG_OH_LINKS_OH5_VFAT16_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT16_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(16).sync_error_cnt;
    regs_read_arr(148)(REG_OH_LINKS_OH5_VFAT16_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT16_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(16).daq_event_cnt;
    regs_read_arr(148)(REG_OH_LINKS_OH5_VFAT16_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT16_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(16).daq_crc_err_cnt;
    regs_read_arr(149)(REG_OH_LINKS_OH5_VFAT17_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(17).sync_good;
    regs_read_arr(149)(REG_OH_LINKS_OH5_VFAT17_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT17_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(17).sync_error_cnt;
    regs_read_arr(149)(REG_OH_LINKS_OH5_VFAT17_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT17_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(17).daq_event_cnt;
    regs_read_arr(149)(REG_OH_LINKS_OH5_VFAT17_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT17_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(17).daq_crc_err_cnt;
    regs_read_arr(150)(REG_OH_LINKS_OH5_VFAT18_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(18).sync_good;
    regs_read_arr(150)(REG_OH_LINKS_OH5_VFAT18_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT18_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(18).sync_error_cnt;
    regs_read_arr(150)(REG_OH_LINKS_OH5_VFAT18_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT18_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(18).daq_event_cnt;
    regs_read_arr(150)(REG_OH_LINKS_OH5_VFAT18_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT18_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(18).daq_crc_err_cnt;
    regs_read_arr(151)(REG_OH_LINKS_OH5_VFAT19_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(19).sync_good;
    regs_read_arr(151)(REG_OH_LINKS_OH5_VFAT19_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT19_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(19).sync_error_cnt;
    regs_read_arr(151)(REG_OH_LINKS_OH5_VFAT19_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT19_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(19).daq_event_cnt;
    regs_read_arr(151)(REG_OH_LINKS_OH5_VFAT19_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT19_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(19).daq_crc_err_cnt;
    regs_read_arr(152)(REG_OH_LINKS_OH5_VFAT20_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(20).sync_good;
    regs_read_arr(152)(REG_OH_LINKS_OH5_VFAT20_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT20_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(20).sync_error_cnt;
    regs_read_arr(152)(REG_OH_LINKS_OH5_VFAT20_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT20_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(20).daq_event_cnt;
    regs_read_arr(152)(REG_OH_LINKS_OH5_VFAT20_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT20_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(20).daq_crc_err_cnt;
    regs_read_arr(153)(REG_OH_LINKS_OH5_VFAT21_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(21).sync_good;
    regs_read_arr(153)(REG_OH_LINKS_OH5_VFAT21_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT21_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(21).sync_error_cnt;
    regs_read_arr(153)(REG_OH_LINKS_OH5_VFAT21_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT21_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(21).daq_event_cnt;
    regs_read_arr(153)(REG_OH_LINKS_OH5_VFAT21_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT21_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(21).daq_crc_err_cnt;
    regs_read_arr(154)(REG_OH_LINKS_OH5_VFAT22_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(22).sync_good;
    regs_read_arr(154)(REG_OH_LINKS_OH5_VFAT22_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT22_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(22).sync_error_cnt;
    regs_read_arr(154)(REG_OH_LINKS_OH5_VFAT22_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT22_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(22).daq_event_cnt;
    regs_read_arr(154)(REG_OH_LINKS_OH5_VFAT22_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT22_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(22).daq_crc_err_cnt;
    regs_read_arr(155)(REG_OH_LINKS_OH5_VFAT23_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(5)(23).sync_good;
    regs_read_arr(155)(REG_OH_LINKS_OH5_VFAT23_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT23_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(5)(23).sync_error_cnt;
    regs_read_arr(155)(REG_OH_LINKS_OH5_VFAT23_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH5_VFAT23_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(5)(23).daq_event_cnt;
    regs_read_arr(155)(REG_OH_LINKS_OH5_VFAT23_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH5_VFAT23_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(5)(23).daq_crc_err_cnt;
    regs_read_arr(156)(REG_OH_LINKS_OH6_GBT0_READY_BIT) <= gbt_link_status_arr_i(6 * g_NUM_GBTS_PER_OH + 0).gbt_rx_ready;
    regs_read_arr(156)(REG_OH_LINKS_OH6_GBT1_READY_BIT) <= gbt_link_status_arr_i(6 * g_NUM_GBTS_PER_OH + 1).gbt_rx_ready;
    regs_read_arr(156)(REG_OH_LINKS_OH6_GBT2_READY_BIT) <= gbt_link_status_arr_i(6 * g_NUM_GBTS_PER_OH + 2).gbt_rx_ready;
    regs_read_arr(156)(REG_OH_LINKS_OH6_GBT0_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(6 * g_NUM_GBTS_PER_OH + 0).gbt_rx_had_not_ready;
    regs_read_arr(156)(REG_OH_LINKS_OH6_GBT1_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(6 * g_NUM_GBTS_PER_OH + 1).gbt_rx_had_not_ready;
    regs_read_arr(156)(REG_OH_LINKS_OH6_GBT2_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(6 * g_NUM_GBTS_PER_OH + 2).gbt_rx_had_not_ready;
    regs_read_arr(156)(REG_OH_LINKS_OH6_GBT0_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(6 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_ovf;
    regs_read_arr(156)(REG_OH_LINKS_OH6_GBT1_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(6 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_ovf;
    regs_read_arr(156)(REG_OH_LINKS_OH6_GBT2_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(6 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_ovf;
    regs_read_arr(156)(REG_OH_LINKS_OH6_GBT0_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(6 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_unf;
    regs_read_arr(156)(REG_OH_LINKS_OH6_GBT1_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(6 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_unf;
    regs_read_arr(156)(REG_OH_LINKS_OH6_GBT2_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(6 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_unf;
    regs_read_arr(157)(REG_OH_LINKS_OH6_VFAT_MASK_MSB downto REG_OH_LINKS_OH6_VFAT_MASK_LSB) <= vfat_mask_arr(6);
    regs_read_arr(158)(REG_OH_LINKS_OH6_VFAT0_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(0).sync_good;
    regs_read_arr(158)(REG_OH_LINKS_OH6_VFAT0_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT0_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(0).sync_error_cnt;
    regs_read_arr(158)(REG_OH_LINKS_OH6_VFAT0_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT0_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(0).daq_event_cnt;
    regs_read_arr(158)(REG_OH_LINKS_OH6_VFAT0_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT0_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(0).daq_crc_err_cnt;
    regs_read_arr(159)(REG_OH_LINKS_OH6_VFAT1_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(1).sync_good;
    regs_read_arr(159)(REG_OH_LINKS_OH6_VFAT1_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT1_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(1).sync_error_cnt;
    regs_read_arr(159)(REG_OH_LINKS_OH6_VFAT1_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT1_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(1).daq_event_cnt;
    regs_read_arr(159)(REG_OH_LINKS_OH6_VFAT1_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT1_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(1).daq_crc_err_cnt;
    regs_read_arr(160)(REG_OH_LINKS_OH6_VFAT2_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(2).sync_good;
    regs_read_arr(160)(REG_OH_LINKS_OH6_VFAT2_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT2_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(2).sync_error_cnt;
    regs_read_arr(160)(REG_OH_LINKS_OH6_VFAT2_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT2_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(2).daq_event_cnt;
    regs_read_arr(160)(REG_OH_LINKS_OH6_VFAT2_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT2_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(2).daq_crc_err_cnt;
    regs_read_arr(161)(REG_OH_LINKS_OH6_VFAT3_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(3).sync_good;
    regs_read_arr(161)(REG_OH_LINKS_OH6_VFAT3_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT3_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(3).sync_error_cnt;
    regs_read_arr(161)(REG_OH_LINKS_OH6_VFAT3_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT3_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(3).daq_event_cnt;
    regs_read_arr(161)(REG_OH_LINKS_OH6_VFAT3_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT3_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(3).daq_crc_err_cnt;
    regs_read_arr(162)(REG_OH_LINKS_OH6_VFAT4_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(4).sync_good;
    regs_read_arr(162)(REG_OH_LINKS_OH6_VFAT4_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT4_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(4).sync_error_cnt;
    regs_read_arr(162)(REG_OH_LINKS_OH6_VFAT4_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT4_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(4).daq_event_cnt;
    regs_read_arr(162)(REG_OH_LINKS_OH6_VFAT4_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT4_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(4).daq_crc_err_cnt;
    regs_read_arr(163)(REG_OH_LINKS_OH6_VFAT5_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(5).sync_good;
    regs_read_arr(163)(REG_OH_LINKS_OH6_VFAT5_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT5_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(5).sync_error_cnt;
    regs_read_arr(163)(REG_OH_LINKS_OH6_VFAT5_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT5_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(5).daq_event_cnt;
    regs_read_arr(163)(REG_OH_LINKS_OH6_VFAT5_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT5_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(5).daq_crc_err_cnt;
    regs_read_arr(164)(REG_OH_LINKS_OH6_VFAT6_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(6).sync_good;
    regs_read_arr(164)(REG_OH_LINKS_OH6_VFAT6_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT6_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(6).sync_error_cnt;
    regs_read_arr(164)(REG_OH_LINKS_OH6_VFAT6_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT6_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(6).daq_event_cnt;
    regs_read_arr(164)(REG_OH_LINKS_OH6_VFAT6_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT6_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(6).daq_crc_err_cnt;
    regs_read_arr(165)(REG_OH_LINKS_OH6_VFAT7_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(7).sync_good;
    regs_read_arr(165)(REG_OH_LINKS_OH6_VFAT7_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT7_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(7).sync_error_cnt;
    regs_read_arr(165)(REG_OH_LINKS_OH6_VFAT7_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT7_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(7).daq_event_cnt;
    regs_read_arr(165)(REG_OH_LINKS_OH6_VFAT7_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT7_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(7).daq_crc_err_cnt;
    regs_read_arr(166)(REG_OH_LINKS_OH6_VFAT8_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(8).sync_good;
    regs_read_arr(166)(REG_OH_LINKS_OH6_VFAT8_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT8_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(8).sync_error_cnt;
    regs_read_arr(166)(REG_OH_LINKS_OH6_VFAT8_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT8_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(8).daq_event_cnt;
    regs_read_arr(166)(REG_OH_LINKS_OH6_VFAT8_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT8_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(8).daq_crc_err_cnt;
    regs_read_arr(167)(REG_OH_LINKS_OH6_VFAT9_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(9).sync_good;
    regs_read_arr(167)(REG_OH_LINKS_OH6_VFAT9_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT9_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(9).sync_error_cnt;
    regs_read_arr(167)(REG_OH_LINKS_OH6_VFAT9_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT9_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(9).daq_event_cnt;
    regs_read_arr(167)(REG_OH_LINKS_OH6_VFAT9_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT9_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(9).daq_crc_err_cnt;
    regs_read_arr(168)(REG_OH_LINKS_OH6_VFAT10_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(10).sync_good;
    regs_read_arr(168)(REG_OH_LINKS_OH6_VFAT10_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT10_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(10).sync_error_cnt;
    regs_read_arr(168)(REG_OH_LINKS_OH6_VFAT10_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT10_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(10).daq_event_cnt;
    regs_read_arr(168)(REG_OH_LINKS_OH6_VFAT10_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT10_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(10).daq_crc_err_cnt;
    regs_read_arr(169)(REG_OH_LINKS_OH6_VFAT11_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(11).sync_good;
    regs_read_arr(169)(REG_OH_LINKS_OH6_VFAT11_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT11_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(11).sync_error_cnt;
    regs_read_arr(169)(REG_OH_LINKS_OH6_VFAT11_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT11_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(11).daq_event_cnt;
    regs_read_arr(169)(REG_OH_LINKS_OH6_VFAT11_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT11_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(11).daq_crc_err_cnt;
    regs_read_arr(170)(REG_OH_LINKS_OH6_VFAT12_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(12).sync_good;
    regs_read_arr(170)(REG_OH_LINKS_OH6_VFAT12_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT12_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(12).sync_error_cnt;
    regs_read_arr(170)(REG_OH_LINKS_OH6_VFAT12_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT12_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(12).daq_event_cnt;
    regs_read_arr(170)(REG_OH_LINKS_OH6_VFAT12_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT12_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(12).daq_crc_err_cnt;
    regs_read_arr(171)(REG_OH_LINKS_OH6_VFAT13_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(13).sync_good;
    regs_read_arr(171)(REG_OH_LINKS_OH6_VFAT13_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT13_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(13).sync_error_cnt;
    regs_read_arr(171)(REG_OH_LINKS_OH6_VFAT13_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT13_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(13).daq_event_cnt;
    regs_read_arr(171)(REG_OH_LINKS_OH6_VFAT13_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT13_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(13).daq_crc_err_cnt;
    regs_read_arr(172)(REG_OH_LINKS_OH6_VFAT14_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(14).sync_good;
    regs_read_arr(172)(REG_OH_LINKS_OH6_VFAT14_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT14_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(14).sync_error_cnt;
    regs_read_arr(172)(REG_OH_LINKS_OH6_VFAT14_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT14_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(14).daq_event_cnt;
    regs_read_arr(172)(REG_OH_LINKS_OH6_VFAT14_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT14_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(14).daq_crc_err_cnt;
    regs_read_arr(173)(REG_OH_LINKS_OH6_VFAT15_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(15).sync_good;
    regs_read_arr(173)(REG_OH_LINKS_OH6_VFAT15_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT15_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(15).sync_error_cnt;
    regs_read_arr(173)(REG_OH_LINKS_OH6_VFAT15_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT15_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(15).daq_event_cnt;
    regs_read_arr(173)(REG_OH_LINKS_OH6_VFAT15_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT15_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(15).daq_crc_err_cnt;
    regs_read_arr(174)(REG_OH_LINKS_OH6_VFAT16_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(16).sync_good;
    regs_read_arr(174)(REG_OH_LINKS_OH6_VFAT16_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT16_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(16).sync_error_cnt;
    regs_read_arr(174)(REG_OH_LINKS_OH6_VFAT16_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT16_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(16).daq_event_cnt;
    regs_read_arr(174)(REG_OH_LINKS_OH6_VFAT16_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT16_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(16).daq_crc_err_cnt;
    regs_read_arr(175)(REG_OH_LINKS_OH6_VFAT17_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(17).sync_good;
    regs_read_arr(175)(REG_OH_LINKS_OH6_VFAT17_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT17_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(17).sync_error_cnt;
    regs_read_arr(175)(REG_OH_LINKS_OH6_VFAT17_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT17_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(17).daq_event_cnt;
    regs_read_arr(175)(REG_OH_LINKS_OH6_VFAT17_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT17_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(17).daq_crc_err_cnt;
    regs_read_arr(176)(REG_OH_LINKS_OH6_VFAT18_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(18).sync_good;
    regs_read_arr(176)(REG_OH_LINKS_OH6_VFAT18_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT18_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(18).sync_error_cnt;
    regs_read_arr(176)(REG_OH_LINKS_OH6_VFAT18_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT18_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(18).daq_event_cnt;
    regs_read_arr(176)(REG_OH_LINKS_OH6_VFAT18_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT18_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(18).daq_crc_err_cnt;
    regs_read_arr(177)(REG_OH_LINKS_OH6_VFAT19_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(19).sync_good;
    regs_read_arr(177)(REG_OH_LINKS_OH6_VFAT19_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT19_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(19).sync_error_cnt;
    regs_read_arr(177)(REG_OH_LINKS_OH6_VFAT19_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT19_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(19).daq_event_cnt;
    regs_read_arr(177)(REG_OH_LINKS_OH6_VFAT19_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT19_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(19).daq_crc_err_cnt;
    regs_read_arr(178)(REG_OH_LINKS_OH6_VFAT20_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(20).sync_good;
    regs_read_arr(178)(REG_OH_LINKS_OH6_VFAT20_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT20_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(20).sync_error_cnt;
    regs_read_arr(178)(REG_OH_LINKS_OH6_VFAT20_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT20_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(20).daq_event_cnt;
    regs_read_arr(178)(REG_OH_LINKS_OH6_VFAT20_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT20_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(20).daq_crc_err_cnt;
    regs_read_arr(179)(REG_OH_LINKS_OH6_VFAT21_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(21).sync_good;
    regs_read_arr(179)(REG_OH_LINKS_OH6_VFAT21_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT21_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(21).sync_error_cnt;
    regs_read_arr(179)(REG_OH_LINKS_OH6_VFAT21_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT21_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(21).daq_event_cnt;
    regs_read_arr(179)(REG_OH_LINKS_OH6_VFAT21_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT21_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(21).daq_crc_err_cnt;
    regs_read_arr(180)(REG_OH_LINKS_OH6_VFAT22_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(22).sync_good;
    regs_read_arr(180)(REG_OH_LINKS_OH6_VFAT22_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT22_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(22).sync_error_cnt;
    regs_read_arr(180)(REG_OH_LINKS_OH6_VFAT22_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT22_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(22).daq_event_cnt;
    regs_read_arr(180)(REG_OH_LINKS_OH6_VFAT22_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT22_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(22).daq_crc_err_cnt;
    regs_read_arr(181)(REG_OH_LINKS_OH6_VFAT23_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(6)(23).sync_good;
    regs_read_arr(181)(REG_OH_LINKS_OH6_VFAT23_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT23_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(6)(23).sync_error_cnt;
    regs_read_arr(181)(REG_OH_LINKS_OH6_VFAT23_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH6_VFAT23_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(6)(23).daq_event_cnt;
    regs_read_arr(181)(REG_OH_LINKS_OH6_VFAT23_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH6_VFAT23_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(6)(23).daq_crc_err_cnt;
    regs_read_arr(182)(REG_OH_LINKS_OH7_GBT0_READY_BIT) <= gbt_link_status_arr_i(7 * g_NUM_GBTS_PER_OH + 0).gbt_rx_ready;
    regs_read_arr(182)(REG_OH_LINKS_OH7_GBT1_READY_BIT) <= gbt_link_status_arr_i(7 * g_NUM_GBTS_PER_OH + 1).gbt_rx_ready;
    regs_read_arr(182)(REG_OH_LINKS_OH7_GBT2_READY_BIT) <= gbt_link_status_arr_i(7 * g_NUM_GBTS_PER_OH + 2).gbt_rx_ready;
    regs_read_arr(182)(REG_OH_LINKS_OH7_GBT0_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(7 * g_NUM_GBTS_PER_OH + 0).gbt_rx_had_not_ready;
    regs_read_arr(182)(REG_OH_LINKS_OH7_GBT1_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(7 * g_NUM_GBTS_PER_OH + 1).gbt_rx_had_not_ready;
    regs_read_arr(182)(REG_OH_LINKS_OH7_GBT2_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(7 * g_NUM_GBTS_PER_OH + 2).gbt_rx_had_not_ready;
    regs_read_arr(182)(REG_OH_LINKS_OH7_GBT0_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(7 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_ovf;
    regs_read_arr(182)(REG_OH_LINKS_OH7_GBT1_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(7 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_ovf;
    regs_read_arr(182)(REG_OH_LINKS_OH7_GBT2_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(7 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_ovf;
    regs_read_arr(182)(REG_OH_LINKS_OH7_GBT0_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(7 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_unf;
    regs_read_arr(182)(REG_OH_LINKS_OH7_GBT1_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(7 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_unf;
    regs_read_arr(182)(REG_OH_LINKS_OH7_GBT2_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(7 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_unf;
    regs_read_arr(183)(REG_OH_LINKS_OH7_VFAT_MASK_MSB downto REG_OH_LINKS_OH7_VFAT_MASK_LSB) <= vfat_mask_arr(7);
    regs_read_arr(184)(REG_OH_LINKS_OH7_VFAT0_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(0).sync_good;
    regs_read_arr(184)(REG_OH_LINKS_OH7_VFAT0_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT0_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(0).sync_error_cnt;
    regs_read_arr(184)(REG_OH_LINKS_OH7_VFAT0_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT0_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(0).daq_event_cnt;
    regs_read_arr(184)(REG_OH_LINKS_OH7_VFAT0_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT0_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(0).daq_crc_err_cnt;
    regs_read_arr(185)(REG_OH_LINKS_OH7_VFAT1_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(1).sync_good;
    regs_read_arr(185)(REG_OH_LINKS_OH7_VFAT1_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT1_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(1).sync_error_cnt;
    regs_read_arr(185)(REG_OH_LINKS_OH7_VFAT1_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT1_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(1).daq_event_cnt;
    regs_read_arr(185)(REG_OH_LINKS_OH7_VFAT1_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT1_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(1).daq_crc_err_cnt;
    regs_read_arr(186)(REG_OH_LINKS_OH7_VFAT2_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(2).sync_good;
    regs_read_arr(186)(REG_OH_LINKS_OH7_VFAT2_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT2_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(2).sync_error_cnt;
    regs_read_arr(186)(REG_OH_LINKS_OH7_VFAT2_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT2_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(2).daq_event_cnt;
    regs_read_arr(186)(REG_OH_LINKS_OH7_VFAT2_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT2_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(2).daq_crc_err_cnt;
    regs_read_arr(187)(REG_OH_LINKS_OH7_VFAT3_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(3).sync_good;
    regs_read_arr(187)(REG_OH_LINKS_OH7_VFAT3_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT3_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(3).sync_error_cnt;
    regs_read_arr(187)(REG_OH_LINKS_OH7_VFAT3_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT3_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(3).daq_event_cnt;
    regs_read_arr(187)(REG_OH_LINKS_OH7_VFAT3_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT3_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(3).daq_crc_err_cnt;
    regs_read_arr(188)(REG_OH_LINKS_OH7_VFAT4_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(4).sync_good;
    regs_read_arr(188)(REG_OH_LINKS_OH7_VFAT4_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT4_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(4).sync_error_cnt;
    regs_read_arr(188)(REG_OH_LINKS_OH7_VFAT4_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT4_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(4).daq_event_cnt;
    regs_read_arr(188)(REG_OH_LINKS_OH7_VFAT4_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT4_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(4).daq_crc_err_cnt;
    regs_read_arr(189)(REG_OH_LINKS_OH7_VFAT5_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(5).sync_good;
    regs_read_arr(189)(REG_OH_LINKS_OH7_VFAT5_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT5_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(5).sync_error_cnt;
    regs_read_arr(189)(REG_OH_LINKS_OH7_VFAT5_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT5_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(5).daq_event_cnt;
    regs_read_arr(189)(REG_OH_LINKS_OH7_VFAT5_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT5_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(5).daq_crc_err_cnt;
    regs_read_arr(190)(REG_OH_LINKS_OH7_VFAT6_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(6).sync_good;
    regs_read_arr(190)(REG_OH_LINKS_OH7_VFAT6_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT6_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(6).sync_error_cnt;
    regs_read_arr(190)(REG_OH_LINKS_OH7_VFAT6_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT6_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(6).daq_event_cnt;
    regs_read_arr(190)(REG_OH_LINKS_OH7_VFAT6_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT6_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(6).daq_crc_err_cnt;
    regs_read_arr(191)(REG_OH_LINKS_OH7_VFAT7_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(7).sync_good;
    regs_read_arr(191)(REG_OH_LINKS_OH7_VFAT7_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT7_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(7).sync_error_cnt;
    regs_read_arr(191)(REG_OH_LINKS_OH7_VFAT7_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT7_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(7).daq_event_cnt;
    regs_read_arr(191)(REG_OH_LINKS_OH7_VFAT7_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT7_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(7).daq_crc_err_cnt;
    regs_read_arr(192)(REG_OH_LINKS_OH7_VFAT8_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(8).sync_good;
    regs_read_arr(192)(REG_OH_LINKS_OH7_VFAT8_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT8_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(8).sync_error_cnt;
    regs_read_arr(192)(REG_OH_LINKS_OH7_VFAT8_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT8_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(8).daq_event_cnt;
    regs_read_arr(192)(REG_OH_LINKS_OH7_VFAT8_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT8_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(8).daq_crc_err_cnt;
    regs_read_arr(193)(REG_OH_LINKS_OH7_VFAT9_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(9).sync_good;
    regs_read_arr(193)(REG_OH_LINKS_OH7_VFAT9_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT9_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(9).sync_error_cnt;
    regs_read_arr(193)(REG_OH_LINKS_OH7_VFAT9_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT9_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(9).daq_event_cnt;
    regs_read_arr(193)(REG_OH_LINKS_OH7_VFAT9_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT9_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(9).daq_crc_err_cnt;
    regs_read_arr(194)(REG_OH_LINKS_OH7_VFAT10_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(10).sync_good;
    regs_read_arr(194)(REG_OH_LINKS_OH7_VFAT10_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT10_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(10).sync_error_cnt;
    regs_read_arr(194)(REG_OH_LINKS_OH7_VFAT10_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT10_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(10).daq_event_cnt;
    regs_read_arr(194)(REG_OH_LINKS_OH7_VFAT10_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT10_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(10).daq_crc_err_cnt;
    regs_read_arr(195)(REG_OH_LINKS_OH7_VFAT11_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(11).sync_good;
    regs_read_arr(195)(REG_OH_LINKS_OH7_VFAT11_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT11_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(11).sync_error_cnt;
    regs_read_arr(195)(REG_OH_LINKS_OH7_VFAT11_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT11_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(11).daq_event_cnt;
    regs_read_arr(195)(REG_OH_LINKS_OH7_VFAT11_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT11_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(11).daq_crc_err_cnt;
    regs_read_arr(196)(REG_OH_LINKS_OH7_VFAT12_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(12).sync_good;
    regs_read_arr(196)(REG_OH_LINKS_OH7_VFAT12_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT12_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(12).sync_error_cnt;
    regs_read_arr(196)(REG_OH_LINKS_OH7_VFAT12_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT12_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(12).daq_event_cnt;
    regs_read_arr(196)(REG_OH_LINKS_OH7_VFAT12_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT12_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(12).daq_crc_err_cnt;
    regs_read_arr(197)(REG_OH_LINKS_OH7_VFAT13_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(13).sync_good;
    regs_read_arr(197)(REG_OH_LINKS_OH7_VFAT13_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT13_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(13).sync_error_cnt;
    regs_read_arr(197)(REG_OH_LINKS_OH7_VFAT13_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT13_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(13).daq_event_cnt;
    regs_read_arr(197)(REG_OH_LINKS_OH7_VFAT13_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT13_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(13).daq_crc_err_cnt;
    regs_read_arr(198)(REG_OH_LINKS_OH7_VFAT14_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(14).sync_good;
    regs_read_arr(198)(REG_OH_LINKS_OH7_VFAT14_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT14_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(14).sync_error_cnt;
    regs_read_arr(198)(REG_OH_LINKS_OH7_VFAT14_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT14_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(14).daq_event_cnt;
    regs_read_arr(198)(REG_OH_LINKS_OH7_VFAT14_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT14_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(14).daq_crc_err_cnt;
    regs_read_arr(199)(REG_OH_LINKS_OH7_VFAT15_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(15).sync_good;
    regs_read_arr(199)(REG_OH_LINKS_OH7_VFAT15_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT15_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(15).sync_error_cnt;
    regs_read_arr(199)(REG_OH_LINKS_OH7_VFAT15_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT15_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(15).daq_event_cnt;
    regs_read_arr(199)(REG_OH_LINKS_OH7_VFAT15_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT15_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(15).daq_crc_err_cnt;
    regs_read_arr(200)(REG_OH_LINKS_OH7_VFAT16_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(16).sync_good;
    regs_read_arr(200)(REG_OH_LINKS_OH7_VFAT16_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT16_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(16).sync_error_cnt;
    regs_read_arr(200)(REG_OH_LINKS_OH7_VFAT16_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT16_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(16).daq_event_cnt;
    regs_read_arr(200)(REG_OH_LINKS_OH7_VFAT16_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT16_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(16).daq_crc_err_cnt;
    regs_read_arr(201)(REG_OH_LINKS_OH7_VFAT17_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(17).sync_good;
    regs_read_arr(201)(REG_OH_LINKS_OH7_VFAT17_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT17_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(17).sync_error_cnt;
    regs_read_arr(201)(REG_OH_LINKS_OH7_VFAT17_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT17_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(17).daq_event_cnt;
    regs_read_arr(201)(REG_OH_LINKS_OH7_VFAT17_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT17_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(17).daq_crc_err_cnt;
    regs_read_arr(202)(REG_OH_LINKS_OH7_VFAT18_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(18).sync_good;
    regs_read_arr(202)(REG_OH_LINKS_OH7_VFAT18_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT18_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(18).sync_error_cnt;
    regs_read_arr(202)(REG_OH_LINKS_OH7_VFAT18_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT18_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(18).daq_event_cnt;
    regs_read_arr(202)(REG_OH_LINKS_OH7_VFAT18_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT18_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(18).daq_crc_err_cnt;
    regs_read_arr(203)(REG_OH_LINKS_OH7_VFAT19_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(19).sync_good;
    regs_read_arr(203)(REG_OH_LINKS_OH7_VFAT19_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT19_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(19).sync_error_cnt;
    regs_read_arr(203)(REG_OH_LINKS_OH7_VFAT19_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT19_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(19).daq_event_cnt;
    regs_read_arr(203)(REG_OH_LINKS_OH7_VFAT19_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT19_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(19).daq_crc_err_cnt;
    regs_read_arr(204)(REG_OH_LINKS_OH7_VFAT20_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(20).sync_good;
    regs_read_arr(204)(REG_OH_LINKS_OH7_VFAT20_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT20_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(20).sync_error_cnt;
    regs_read_arr(204)(REG_OH_LINKS_OH7_VFAT20_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT20_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(20).daq_event_cnt;
    regs_read_arr(204)(REG_OH_LINKS_OH7_VFAT20_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT20_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(20).daq_crc_err_cnt;
    regs_read_arr(205)(REG_OH_LINKS_OH7_VFAT21_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(21).sync_good;
    regs_read_arr(205)(REG_OH_LINKS_OH7_VFAT21_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT21_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(21).sync_error_cnt;
    regs_read_arr(205)(REG_OH_LINKS_OH7_VFAT21_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT21_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(21).daq_event_cnt;
    regs_read_arr(205)(REG_OH_LINKS_OH7_VFAT21_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT21_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(21).daq_crc_err_cnt;
    regs_read_arr(206)(REG_OH_LINKS_OH7_VFAT22_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(22).sync_good;
    regs_read_arr(206)(REG_OH_LINKS_OH7_VFAT22_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT22_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(22).sync_error_cnt;
    regs_read_arr(206)(REG_OH_LINKS_OH7_VFAT22_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT22_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(22).daq_event_cnt;
    regs_read_arr(206)(REG_OH_LINKS_OH7_VFAT22_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT22_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(22).daq_crc_err_cnt;
    regs_read_arr(207)(REG_OH_LINKS_OH7_VFAT23_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(7)(23).sync_good;
    regs_read_arr(207)(REG_OH_LINKS_OH7_VFAT23_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT23_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(7)(23).sync_error_cnt;
    regs_read_arr(207)(REG_OH_LINKS_OH7_VFAT23_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH7_VFAT23_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(7)(23).daq_event_cnt;
    regs_read_arr(207)(REG_OH_LINKS_OH7_VFAT23_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH7_VFAT23_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(7)(23).daq_crc_err_cnt;
    regs_read_arr(208)(REG_OH_LINKS_OH8_GBT0_READY_BIT) <= gbt_link_status_arr_i(8 * g_NUM_GBTS_PER_OH + 0).gbt_rx_ready;
    regs_read_arr(208)(REG_OH_LINKS_OH8_GBT1_READY_BIT) <= gbt_link_status_arr_i(8 * g_NUM_GBTS_PER_OH + 1).gbt_rx_ready;
    regs_read_arr(208)(REG_OH_LINKS_OH8_GBT2_READY_BIT) <= gbt_link_status_arr_i(8 * g_NUM_GBTS_PER_OH + 2).gbt_rx_ready;
    regs_read_arr(208)(REG_OH_LINKS_OH8_GBT0_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(8 * g_NUM_GBTS_PER_OH + 0).gbt_rx_had_not_ready;
    regs_read_arr(208)(REG_OH_LINKS_OH8_GBT1_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(8 * g_NUM_GBTS_PER_OH + 1).gbt_rx_had_not_ready;
    regs_read_arr(208)(REG_OH_LINKS_OH8_GBT2_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(8 * g_NUM_GBTS_PER_OH + 2).gbt_rx_had_not_ready;
    regs_read_arr(208)(REG_OH_LINKS_OH8_GBT0_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(8 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_ovf;
    regs_read_arr(208)(REG_OH_LINKS_OH8_GBT1_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(8 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_ovf;
    regs_read_arr(208)(REG_OH_LINKS_OH8_GBT2_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(8 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_ovf;
    regs_read_arr(208)(REG_OH_LINKS_OH8_GBT0_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(8 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_unf;
    regs_read_arr(208)(REG_OH_LINKS_OH8_GBT1_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(8 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_unf;
    regs_read_arr(208)(REG_OH_LINKS_OH8_GBT2_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(8 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_unf;
    regs_read_arr(209)(REG_OH_LINKS_OH8_VFAT_MASK_MSB downto REG_OH_LINKS_OH8_VFAT_MASK_LSB) <= vfat_mask_arr(8);
    regs_read_arr(210)(REG_OH_LINKS_OH8_VFAT0_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(0).sync_good;
    regs_read_arr(210)(REG_OH_LINKS_OH8_VFAT0_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT0_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(0).sync_error_cnt;
    regs_read_arr(210)(REG_OH_LINKS_OH8_VFAT0_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT0_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(0).daq_event_cnt;
    regs_read_arr(210)(REG_OH_LINKS_OH8_VFAT0_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT0_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(0).daq_crc_err_cnt;
    regs_read_arr(211)(REG_OH_LINKS_OH8_VFAT1_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(1).sync_good;
    regs_read_arr(211)(REG_OH_LINKS_OH8_VFAT1_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT1_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(1).sync_error_cnt;
    regs_read_arr(211)(REG_OH_LINKS_OH8_VFAT1_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT1_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(1).daq_event_cnt;
    regs_read_arr(211)(REG_OH_LINKS_OH8_VFAT1_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT1_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(1).daq_crc_err_cnt;
    regs_read_arr(212)(REG_OH_LINKS_OH8_VFAT2_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(2).sync_good;
    regs_read_arr(212)(REG_OH_LINKS_OH8_VFAT2_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT2_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(2).sync_error_cnt;
    regs_read_arr(212)(REG_OH_LINKS_OH8_VFAT2_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT2_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(2).daq_event_cnt;
    regs_read_arr(212)(REG_OH_LINKS_OH8_VFAT2_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT2_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(2).daq_crc_err_cnt;
    regs_read_arr(213)(REG_OH_LINKS_OH8_VFAT3_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(3).sync_good;
    regs_read_arr(213)(REG_OH_LINKS_OH8_VFAT3_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT3_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(3).sync_error_cnt;
    regs_read_arr(213)(REG_OH_LINKS_OH8_VFAT3_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT3_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(3).daq_event_cnt;
    regs_read_arr(213)(REG_OH_LINKS_OH8_VFAT3_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT3_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(3).daq_crc_err_cnt;
    regs_read_arr(214)(REG_OH_LINKS_OH8_VFAT4_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(4).sync_good;
    regs_read_arr(214)(REG_OH_LINKS_OH8_VFAT4_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT4_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(4).sync_error_cnt;
    regs_read_arr(214)(REG_OH_LINKS_OH8_VFAT4_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT4_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(4).daq_event_cnt;
    regs_read_arr(214)(REG_OH_LINKS_OH8_VFAT4_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT4_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(4).daq_crc_err_cnt;
    regs_read_arr(215)(REG_OH_LINKS_OH8_VFAT5_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(5).sync_good;
    regs_read_arr(215)(REG_OH_LINKS_OH8_VFAT5_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT5_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(5).sync_error_cnt;
    regs_read_arr(215)(REG_OH_LINKS_OH8_VFAT5_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT5_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(5).daq_event_cnt;
    regs_read_arr(215)(REG_OH_LINKS_OH8_VFAT5_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT5_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(5).daq_crc_err_cnt;
    regs_read_arr(216)(REG_OH_LINKS_OH8_VFAT6_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(6).sync_good;
    regs_read_arr(216)(REG_OH_LINKS_OH8_VFAT6_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT6_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(6).sync_error_cnt;
    regs_read_arr(216)(REG_OH_LINKS_OH8_VFAT6_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT6_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(6).daq_event_cnt;
    regs_read_arr(216)(REG_OH_LINKS_OH8_VFAT6_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT6_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(6).daq_crc_err_cnt;
    regs_read_arr(217)(REG_OH_LINKS_OH8_VFAT7_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(7).sync_good;
    regs_read_arr(217)(REG_OH_LINKS_OH8_VFAT7_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT7_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(7).sync_error_cnt;
    regs_read_arr(217)(REG_OH_LINKS_OH8_VFAT7_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT7_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(7).daq_event_cnt;
    regs_read_arr(217)(REG_OH_LINKS_OH8_VFAT7_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT7_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(7).daq_crc_err_cnt;
    regs_read_arr(218)(REG_OH_LINKS_OH8_VFAT8_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(8).sync_good;
    regs_read_arr(218)(REG_OH_LINKS_OH8_VFAT8_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT8_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(8).sync_error_cnt;
    regs_read_arr(218)(REG_OH_LINKS_OH8_VFAT8_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT8_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(8).daq_event_cnt;
    regs_read_arr(218)(REG_OH_LINKS_OH8_VFAT8_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT8_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(8).daq_crc_err_cnt;
    regs_read_arr(219)(REG_OH_LINKS_OH8_VFAT9_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(9).sync_good;
    regs_read_arr(219)(REG_OH_LINKS_OH8_VFAT9_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT9_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(9).sync_error_cnt;
    regs_read_arr(219)(REG_OH_LINKS_OH8_VFAT9_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT9_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(9).daq_event_cnt;
    regs_read_arr(219)(REG_OH_LINKS_OH8_VFAT9_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT9_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(9).daq_crc_err_cnt;
    regs_read_arr(220)(REG_OH_LINKS_OH8_VFAT10_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(10).sync_good;
    regs_read_arr(220)(REG_OH_LINKS_OH8_VFAT10_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT10_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(10).sync_error_cnt;
    regs_read_arr(220)(REG_OH_LINKS_OH8_VFAT10_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT10_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(10).daq_event_cnt;
    regs_read_arr(220)(REG_OH_LINKS_OH8_VFAT10_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT10_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(10).daq_crc_err_cnt;
    regs_read_arr(221)(REG_OH_LINKS_OH8_VFAT11_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(11).sync_good;
    regs_read_arr(221)(REG_OH_LINKS_OH8_VFAT11_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT11_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(11).sync_error_cnt;
    regs_read_arr(221)(REG_OH_LINKS_OH8_VFAT11_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT11_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(11).daq_event_cnt;
    regs_read_arr(221)(REG_OH_LINKS_OH8_VFAT11_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT11_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(11).daq_crc_err_cnt;
    regs_read_arr(222)(REG_OH_LINKS_OH8_VFAT12_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(12).sync_good;
    regs_read_arr(222)(REG_OH_LINKS_OH8_VFAT12_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT12_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(12).sync_error_cnt;
    regs_read_arr(222)(REG_OH_LINKS_OH8_VFAT12_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT12_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(12).daq_event_cnt;
    regs_read_arr(222)(REG_OH_LINKS_OH8_VFAT12_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT12_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(12).daq_crc_err_cnt;
    regs_read_arr(223)(REG_OH_LINKS_OH8_VFAT13_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(13).sync_good;
    regs_read_arr(223)(REG_OH_LINKS_OH8_VFAT13_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT13_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(13).sync_error_cnt;
    regs_read_arr(223)(REG_OH_LINKS_OH8_VFAT13_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT13_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(13).daq_event_cnt;
    regs_read_arr(223)(REG_OH_LINKS_OH8_VFAT13_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT13_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(13).daq_crc_err_cnt;
    regs_read_arr(224)(REG_OH_LINKS_OH8_VFAT14_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(14).sync_good;
    regs_read_arr(224)(REG_OH_LINKS_OH8_VFAT14_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT14_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(14).sync_error_cnt;
    regs_read_arr(224)(REG_OH_LINKS_OH8_VFAT14_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT14_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(14).daq_event_cnt;
    regs_read_arr(224)(REG_OH_LINKS_OH8_VFAT14_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT14_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(14).daq_crc_err_cnt;
    regs_read_arr(225)(REG_OH_LINKS_OH8_VFAT15_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(15).sync_good;
    regs_read_arr(225)(REG_OH_LINKS_OH8_VFAT15_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT15_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(15).sync_error_cnt;
    regs_read_arr(225)(REG_OH_LINKS_OH8_VFAT15_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT15_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(15).daq_event_cnt;
    regs_read_arr(225)(REG_OH_LINKS_OH8_VFAT15_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT15_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(15).daq_crc_err_cnt;
    regs_read_arr(226)(REG_OH_LINKS_OH8_VFAT16_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(16).sync_good;
    regs_read_arr(226)(REG_OH_LINKS_OH8_VFAT16_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT16_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(16).sync_error_cnt;
    regs_read_arr(226)(REG_OH_LINKS_OH8_VFAT16_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT16_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(16).daq_event_cnt;
    regs_read_arr(226)(REG_OH_LINKS_OH8_VFAT16_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT16_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(16).daq_crc_err_cnt;
    regs_read_arr(227)(REG_OH_LINKS_OH8_VFAT17_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(17).sync_good;
    regs_read_arr(227)(REG_OH_LINKS_OH8_VFAT17_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT17_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(17).sync_error_cnt;
    regs_read_arr(227)(REG_OH_LINKS_OH8_VFAT17_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT17_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(17).daq_event_cnt;
    regs_read_arr(227)(REG_OH_LINKS_OH8_VFAT17_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT17_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(17).daq_crc_err_cnt;
    regs_read_arr(228)(REG_OH_LINKS_OH8_VFAT18_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(18).sync_good;
    regs_read_arr(228)(REG_OH_LINKS_OH8_VFAT18_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT18_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(18).sync_error_cnt;
    regs_read_arr(228)(REG_OH_LINKS_OH8_VFAT18_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT18_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(18).daq_event_cnt;
    regs_read_arr(228)(REG_OH_LINKS_OH8_VFAT18_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT18_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(18).daq_crc_err_cnt;
    regs_read_arr(229)(REG_OH_LINKS_OH8_VFAT19_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(19).sync_good;
    regs_read_arr(229)(REG_OH_LINKS_OH8_VFAT19_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT19_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(19).sync_error_cnt;
    regs_read_arr(229)(REG_OH_LINKS_OH8_VFAT19_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT19_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(19).daq_event_cnt;
    regs_read_arr(229)(REG_OH_LINKS_OH8_VFAT19_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT19_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(19).daq_crc_err_cnt;
    regs_read_arr(230)(REG_OH_LINKS_OH8_VFAT20_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(20).sync_good;
    regs_read_arr(230)(REG_OH_LINKS_OH8_VFAT20_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT20_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(20).sync_error_cnt;
    regs_read_arr(230)(REG_OH_LINKS_OH8_VFAT20_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT20_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(20).daq_event_cnt;
    regs_read_arr(230)(REG_OH_LINKS_OH8_VFAT20_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT20_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(20).daq_crc_err_cnt;
    regs_read_arr(231)(REG_OH_LINKS_OH8_VFAT21_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(21).sync_good;
    regs_read_arr(231)(REG_OH_LINKS_OH8_VFAT21_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT21_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(21).sync_error_cnt;
    regs_read_arr(231)(REG_OH_LINKS_OH8_VFAT21_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT21_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(21).daq_event_cnt;
    regs_read_arr(231)(REG_OH_LINKS_OH8_VFAT21_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT21_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(21).daq_crc_err_cnt;
    regs_read_arr(232)(REG_OH_LINKS_OH8_VFAT22_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(22).sync_good;
    regs_read_arr(232)(REG_OH_LINKS_OH8_VFAT22_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT22_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(22).sync_error_cnt;
    regs_read_arr(232)(REG_OH_LINKS_OH8_VFAT22_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT22_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(22).daq_event_cnt;
    regs_read_arr(232)(REG_OH_LINKS_OH8_VFAT22_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT22_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(22).daq_crc_err_cnt;
    regs_read_arr(233)(REG_OH_LINKS_OH8_VFAT23_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(8)(23).sync_good;
    regs_read_arr(233)(REG_OH_LINKS_OH8_VFAT23_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT23_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(8)(23).sync_error_cnt;
    regs_read_arr(233)(REG_OH_LINKS_OH8_VFAT23_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH8_VFAT23_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(8)(23).daq_event_cnt;
    regs_read_arr(233)(REG_OH_LINKS_OH8_VFAT23_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH8_VFAT23_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(8)(23).daq_crc_err_cnt;
    regs_read_arr(234)(REG_OH_LINKS_OH9_GBT0_READY_BIT) <= gbt_link_status_arr_i(9 * g_NUM_GBTS_PER_OH + 0).gbt_rx_ready;
    regs_read_arr(234)(REG_OH_LINKS_OH9_GBT1_READY_BIT) <= gbt_link_status_arr_i(9 * g_NUM_GBTS_PER_OH + 1).gbt_rx_ready;
    regs_read_arr(234)(REG_OH_LINKS_OH9_GBT2_READY_BIT) <= gbt_link_status_arr_i(9 * g_NUM_GBTS_PER_OH + 2).gbt_rx_ready;
    regs_read_arr(234)(REG_OH_LINKS_OH9_GBT0_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(9 * g_NUM_GBTS_PER_OH + 0).gbt_rx_had_not_ready;
    regs_read_arr(234)(REG_OH_LINKS_OH9_GBT1_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(9 * g_NUM_GBTS_PER_OH + 1).gbt_rx_had_not_ready;
    regs_read_arr(234)(REG_OH_LINKS_OH9_GBT2_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(9 * g_NUM_GBTS_PER_OH + 2).gbt_rx_had_not_ready;
    regs_read_arr(234)(REG_OH_LINKS_OH9_GBT0_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(9 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_ovf;
    regs_read_arr(234)(REG_OH_LINKS_OH9_GBT1_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(9 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_ovf;
    regs_read_arr(234)(REG_OH_LINKS_OH9_GBT2_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(9 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_ovf;
    regs_read_arr(234)(REG_OH_LINKS_OH9_GBT0_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(9 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_unf;
    regs_read_arr(234)(REG_OH_LINKS_OH9_GBT1_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(9 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_unf;
    regs_read_arr(234)(REG_OH_LINKS_OH9_GBT2_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(9 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_unf;
    regs_read_arr(235)(REG_OH_LINKS_OH9_VFAT_MASK_MSB downto REG_OH_LINKS_OH9_VFAT_MASK_LSB) <= vfat_mask_arr(9);
    regs_read_arr(236)(REG_OH_LINKS_OH9_VFAT0_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(0).sync_good;
    regs_read_arr(236)(REG_OH_LINKS_OH9_VFAT0_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT0_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(0).sync_error_cnt;
    regs_read_arr(236)(REG_OH_LINKS_OH9_VFAT0_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT0_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(0).daq_event_cnt;
    regs_read_arr(236)(REG_OH_LINKS_OH9_VFAT0_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT0_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(0).daq_crc_err_cnt;
    regs_read_arr(237)(REG_OH_LINKS_OH9_VFAT1_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(1).sync_good;
    regs_read_arr(237)(REG_OH_LINKS_OH9_VFAT1_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT1_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(1).sync_error_cnt;
    regs_read_arr(237)(REG_OH_LINKS_OH9_VFAT1_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT1_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(1).daq_event_cnt;
    regs_read_arr(237)(REG_OH_LINKS_OH9_VFAT1_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT1_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(1).daq_crc_err_cnt;
    regs_read_arr(238)(REG_OH_LINKS_OH9_VFAT2_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(2).sync_good;
    regs_read_arr(238)(REG_OH_LINKS_OH9_VFAT2_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT2_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(2).sync_error_cnt;
    regs_read_arr(238)(REG_OH_LINKS_OH9_VFAT2_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT2_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(2).daq_event_cnt;
    regs_read_arr(238)(REG_OH_LINKS_OH9_VFAT2_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT2_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(2).daq_crc_err_cnt;
    regs_read_arr(239)(REG_OH_LINKS_OH9_VFAT3_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(3).sync_good;
    regs_read_arr(239)(REG_OH_LINKS_OH9_VFAT3_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT3_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(3).sync_error_cnt;
    regs_read_arr(239)(REG_OH_LINKS_OH9_VFAT3_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT3_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(3).daq_event_cnt;
    regs_read_arr(239)(REG_OH_LINKS_OH9_VFAT3_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT3_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(3).daq_crc_err_cnt;
    regs_read_arr(240)(REG_OH_LINKS_OH9_VFAT4_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(4).sync_good;
    regs_read_arr(240)(REG_OH_LINKS_OH9_VFAT4_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT4_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(4).sync_error_cnt;
    regs_read_arr(240)(REG_OH_LINKS_OH9_VFAT4_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT4_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(4).daq_event_cnt;
    regs_read_arr(240)(REG_OH_LINKS_OH9_VFAT4_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT4_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(4).daq_crc_err_cnt;
    regs_read_arr(241)(REG_OH_LINKS_OH9_VFAT5_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(5).sync_good;
    regs_read_arr(241)(REG_OH_LINKS_OH9_VFAT5_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT5_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(5).sync_error_cnt;
    regs_read_arr(241)(REG_OH_LINKS_OH9_VFAT5_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT5_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(5).daq_event_cnt;
    regs_read_arr(241)(REG_OH_LINKS_OH9_VFAT5_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT5_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(5).daq_crc_err_cnt;
    regs_read_arr(242)(REG_OH_LINKS_OH9_VFAT6_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(6).sync_good;
    regs_read_arr(242)(REG_OH_LINKS_OH9_VFAT6_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT6_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(6).sync_error_cnt;
    regs_read_arr(242)(REG_OH_LINKS_OH9_VFAT6_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT6_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(6).daq_event_cnt;
    regs_read_arr(242)(REG_OH_LINKS_OH9_VFAT6_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT6_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(6).daq_crc_err_cnt;
    regs_read_arr(243)(REG_OH_LINKS_OH9_VFAT7_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(7).sync_good;
    regs_read_arr(243)(REG_OH_LINKS_OH9_VFAT7_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT7_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(7).sync_error_cnt;
    regs_read_arr(243)(REG_OH_LINKS_OH9_VFAT7_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT7_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(7).daq_event_cnt;
    regs_read_arr(243)(REG_OH_LINKS_OH9_VFAT7_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT7_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(7).daq_crc_err_cnt;
    regs_read_arr(244)(REG_OH_LINKS_OH9_VFAT8_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(8).sync_good;
    regs_read_arr(244)(REG_OH_LINKS_OH9_VFAT8_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT8_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(8).sync_error_cnt;
    regs_read_arr(244)(REG_OH_LINKS_OH9_VFAT8_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT8_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(8).daq_event_cnt;
    regs_read_arr(244)(REG_OH_LINKS_OH9_VFAT8_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT8_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(8).daq_crc_err_cnt;
    regs_read_arr(245)(REG_OH_LINKS_OH9_VFAT9_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(9).sync_good;
    regs_read_arr(245)(REG_OH_LINKS_OH9_VFAT9_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT9_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(9).sync_error_cnt;
    regs_read_arr(245)(REG_OH_LINKS_OH9_VFAT9_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT9_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(9).daq_event_cnt;
    regs_read_arr(245)(REG_OH_LINKS_OH9_VFAT9_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT9_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(9).daq_crc_err_cnt;
    regs_read_arr(246)(REG_OH_LINKS_OH9_VFAT10_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(10).sync_good;
    regs_read_arr(246)(REG_OH_LINKS_OH9_VFAT10_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT10_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(10).sync_error_cnt;
    regs_read_arr(246)(REG_OH_LINKS_OH9_VFAT10_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT10_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(10).daq_event_cnt;
    regs_read_arr(246)(REG_OH_LINKS_OH9_VFAT10_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT10_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(10).daq_crc_err_cnt;
    regs_read_arr(247)(REG_OH_LINKS_OH9_VFAT11_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(11).sync_good;
    regs_read_arr(247)(REG_OH_LINKS_OH9_VFAT11_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT11_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(11).sync_error_cnt;
    regs_read_arr(247)(REG_OH_LINKS_OH9_VFAT11_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT11_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(11).daq_event_cnt;
    regs_read_arr(247)(REG_OH_LINKS_OH9_VFAT11_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT11_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(11).daq_crc_err_cnt;
    regs_read_arr(248)(REG_OH_LINKS_OH9_VFAT12_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(12).sync_good;
    regs_read_arr(248)(REG_OH_LINKS_OH9_VFAT12_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT12_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(12).sync_error_cnt;
    regs_read_arr(248)(REG_OH_LINKS_OH9_VFAT12_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT12_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(12).daq_event_cnt;
    regs_read_arr(248)(REG_OH_LINKS_OH9_VFAT12_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT12_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(12).daq_crc_err_cnt;
    regs_read_arr(249)(REG_OH_LINKS_OH9_VFAT13_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(13).sync_good;
    regs_read_arr(249)(REG_OH_LINKS_OH9_VFAT13_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT13_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(13).sync_error_cnt;
    regs_read_arr(249)(REG_OH_LINKS_OH9_VFAT13_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT13_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(13).daq_event_cnt;
    regs_read_arr(249)(REG_OH_LINKS_OH9_VFAT13_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT13_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(13).daq_crc_err_cnt;
    regs_read_arr(250)(REG_OH_LINKS_OH9_VFAT14_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(14).sync_good;
    regs_read_arr(250)(REG_OH_LINKS_OH9_VFAT14_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT14_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(14).sync_error_cnt;
    regs_read_arr(250)(REG_OH_LINKS_OH9_VFAT14_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT14_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(14).daq_event_cnt;
    regs_read_arr(250)(REG_OH_LINKS_OH9_VFAT14_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT14_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(14).daq_crc_err_cnt;
    regs_read_arr(251)(REG_OH_LINKS_OH9_VFAT15_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(15).sync_good;
    regs_read_arr(251)(REG_OH_LINKS_OH9_VFAT15_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT15_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(15).sync_error_cnt;
    regs_read_arr(251)(REG_OH_LINKS_OH9_VFAT15_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT15_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(15).daq_event_cnt;
    regs_read_arr(251)(REG_OH_LINKS_OH9_VFAT15_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT15_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(15).daq_crc_err_cnt;
    regs_read_arr(252)(REG_OH_LINKS_OH9_VFAT16_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(16).sync_good;
    regs_read_arr(252)(REG_OH_LINKS_OH9_VFAT16_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT16_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(16).sync_error_cnt;
    regs_read_arr(252)(REG_OH_LINKS_OH9_VFAT16_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT16_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(16).daq_event_cnt;
    regs_read_arr(252)(REG_OH_LINKS_OH9_VFAT16_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT16_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(16).daq_crc_err_cnt;
    regs_read_arr(253)(REG_OH_LINKS_OH9_VFAT17_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(17).sync_good;
    regs_read_arr(253)(REG_OH_LINKS_OH9_VFAT17_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT17_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(17).sync_error_cnt;
    regs_read_arr(253)(REG_OH_LINKS_OH9_VFAT17_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT17_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(17).daq_event_cnt;
    regs_read_arr(253)(REG_OH_LINKS_OH9_VFAT17_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT17_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(17).daq_crc_err_cnt;
    regs_read_arr(254)(REG_OH_LINKS_OH9_VFAT18_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(18).sync_good;
    regs_read_arr(254)(REG_OH_LINKS_OH9_VFAT18_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT18_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(18).sync_error_cnt;
    regs_read_arr(254)(REG_OH_LINKS_OH9_VFAT18_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT18_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(18).daq_event_cnt;
    regs_read_arr(254)(REG_OH_LINKS_OH9_VFAT18_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT18_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(18).daq_crc_err_cnt;
    regs_read_arr(255)(REG_OH_LINKS_OH9_VFAT19_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(19).sync_good;
    regs_read_arr(255)(REG_OH_LINKS_OH9_VFAT19_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT19_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(19).sync_error_cnt;
    regs_read_arr(255)(REG_OH_LINKS_OH9_VFAT19_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT19_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(19).daq_event_cnt;
    regs_read_arr(255)(REG_OH_LINKS_OH9_VFAT19_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT19_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(19).daq_crc_err_cnt;
    regs_read_arr(256)(REG_OH_LINKS_OH9_VFAT20_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(20).sync_good;
    regs_read_arr(256)(REG_OH_LINKS_OH9_VFAT20_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT20_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(20).sync_error_cnt;
    regs_read_arr(256)(REG_OH_LINKS_OH9_VFAT20_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT20_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(20).daq_event_cnt;
    regs_read_arr(256)(REG_OH_LINKS_OH9_VFAT20_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT20_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(20).daq_crc_err_cnt;
    regs_read_arr(257)(REG_OH_LINKS_OH9_VFAT21_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(21).sync_good;
    regs_read_arr(257)(REG_OH_LINKS_OH9_VFAT21_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT21_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(21).sync_error_cnt;
    regs_read_arr(257)(REG_OH_LINKS_OH9_VFAT21_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT21_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(21).daq_event_cnt;
    regs_read_arr(257)(REG_OH_LINKS_OH9_VFAT21_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT21_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(21).daq_crc_err_cnt;
    regs_read_arr(258)(REG_OH_LINKS_OH9_VFAT22_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(22).sync_good;
    regs_read_arr(258)(REG_OH_LINKS_OH9_VFAT22_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT22_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(22).sync_error_cnt;
    regs_read_arr(258)(REG_OH_LINKS_OH9_VFAT22_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT22_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(22).daq_event_cnt;
    regs_read_arr(258)(REG_OH_LINKS_OH9_VFAT22_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT22_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(22).daq_crc_err_cnt;
    regs_read_arr(259)(REG_OH_LINKS_OH9_VFAT23_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(9)(23).sync_good;
    regs_read_arr(259)(REG_OH_LINKS_OH9_VFAT23_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT23_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(9)(23).sync_error_cnt;
    regs_read_arr(259)(REG_OH_LINKS_OH9_VFAT23_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH9_VFAT23_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(9)(23).daq_event_cnt;
    regs_read_arr(259)(REG_OH_LINKS_OH9_VFAT23_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH9_VFAT23_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(9)(23).daq_crc_err_cnt;
    regs_read_arr(260)(REG_OH_LINKS_OH10_GBT0_READY_BIT) <= gbt_link_status_arr_i(10 * g_NUM_GBTS_PER_OH + 0).gbt_rx_ready;
    regs_read_arr(260)(REG_OH_LINKS_OH10_GBT1_READY_BIT) <= gbt_link_status_arr_i(10 * g_NUM_GBTS_PER_OH + 1).gbt_rx_ready;
    regs_read_arr(260)(REG_OH_LINKS_OH10_GBT2_READY_BIT) <= gbt_link_status_arr_i(10 * g_NUM_GBTS_PER_OH + 2).gbt_rx_ready;
    regs_read_arr(260)(REG_OH_LINKS_OH10_GBT0_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(10 * g_NUM_GBTS_PER_OH + 0).gbt_rx_had_not_ready;
    regs_read_arr(260)(REG_OH_LINKS_OH10_GBT1_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(10 * g_NUM_GBTS_PER_OH + 1).gbt_rx_had_not_ready;
    regs_read_arr(260)(REG_OH_LINKS_OH10_GBT2_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(10 * g_NUM_GBTS_PER_OH + 2).gbt_rx_had_not_ready;
    regs_read_arr(260)(REG_OH_LINKS_OH10_GBT0_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(10 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_ovf;
    regs_read_arr(260)(REG_OH_LINKS_OH10_GBT1_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(10 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_ovf;
    regs_read_arr(260)(REG_OH_LINKS_OH10_GBT2_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(10 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_ovf;
    regs_read_arr(260)(REG_OH_LINKS_OH10_GBT0_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(10 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_unf;
    regs_read_arr(260)(REG_OH_LINKS_OH10_GBT1_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(10 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_unf;
    regs_read_arr(260)(REG_OH_LINKS_OH10_GBT2_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(10 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_unf;
    regs_read_arr(261)(REG_OH_LINKS_OH10_VFAT_MASK_MSB downto REG_OH_LINKS_OH10_VFAT_MASK_LSB) <= vfat_mask_arr(10);
    regs_read_arr(262)(REG_OH_LINKS_OH10_VFAT0_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(0).sync_good;
    regs_read_arr(262)(REG_OH_LINKS_OH10_VFAT0_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT0_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(0).sync_error_cnt;
    regs_read_arr(262)(REG_OH_LINKS_OH10_VFAT0_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT0_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(0).daq_event_cnt;
    regs_read_arr(262)(REG_OH_LINKS_OH10_VFAT0_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT0_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(0).daq_crc_err_cnt;
    regs_read_arr(263)(REG_OH_LINKS_OH10_VFAT1_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(1).sync_good;
    regs_read_arr(263)(REG_OH_LINKS_OH10_VFAT1_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT1_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(1).sync_error_cnt;
    regs_read_arr(263)(REG_OH_LINKS_OH10_VFAT1_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT1_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(1).daq_event_cnt;
    regs_read_arr(263)(REG_OH_LINKS_OH10_VFAT1_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT1_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(1).daq_crc_err_cnt;
    regs_read_arr(264)(REG_OH_LINKS_OH10_VFAT2_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(2).sync_good;
    regs_read_arr(264)(REG_OH_LINKS_OH10_VFAT2_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT2_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(2).sync_error_cnt;
    regs_read_arr(264)(REG_OH_LINKS_OH10_VFAT2_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT2_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(2).daq_event_cnt;
    regs_read_arr(264)(REG_OH_LINKS_OH10_VFAT2_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT2_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(2).daq_crc_err_cnt;
    regs_read_arr(265)(REG_OH_LINKS_OH10_VFAT3_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(3).sync_good;
    regs_read_arr(265)(REG_OH_LINKS_OH10_VFAT3_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT3_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(3).sync_error_cnt;
    regs_read_arr(265)(REG_OH_LINKS_OH10_VFAT3_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT3_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(3).daq_event_cnt;
    regs_read_arr(265)(REG_OH_LINKS_OH10_VFAT3_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT3_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(3).daq_crc_err_cnt;
    regs_read_arr(266)(REG_OH_LINKS_OH10_VFAT4_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(4).sync_good;
    regs_read_arr(266)(REG_OH_LINKS_OH10_VFAT4_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT4_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(4).sync_error_cnt;
    regs_read_arr(266)(REG_OH_LINKS_OH10_VFAT4_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT4_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(4).daq_event_cnt;
    regs_read_arr(266)(REG_OH_LINKS_OH10_VFAT4_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT4_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(4).daq_crc_err_cnt;
    regs_read_arr(267)(REG_OH_LINKS_OH10_VFAT5_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(5).sync_good;
    regs_read_arr(267)(REG_OH_LINKS_OH10_VFAT5_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT5_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(5).sync_error_cnt;
    regs_read_arr(267)(REG_OH_LINKS_OH10_VFAT5_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT5_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(5).daq_event_cnt;
    regs_read_arr(267)(REG_OH_LINKS_OH10_VFAT5_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT5_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(5).daq_crc_err_cnt;
    regs_read_arr(268)(REG_OH_LINKS_OH10_VFAT6_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(6).sync_good;
    regs_read_arr(268)(REG_OH_LINKS_OH10_VFAT6_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT6_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(6).sync_error_cnt;
    regs_read_arr(268)(REG_OH_LINKS_OH10_VFAT6_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT6_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(6).daq_event_cnt;
    regs_read_arr(268)(REG_OH_LINKS_OH10_VFAT6_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT6_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(6).daq_crc_err_cnt;
    regs_read_arr(269)(REG_OH_LINKS_OH10_VFAT7_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(7).sync_good;
    regs_read_arr(269)(REG_OH_LINKS_OH10_VFAT7_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT7_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(7).sync_error_cnt;
    regs_read_arr(269)(REG_OH_LINKS_OH10_VFAT7_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT7_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(7).daq_event_cnt;
    regs_read_arr(269)(REG_OH_LINKS_OH10_VFAT7_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT7_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(7).daq_crc_err_cnt;
    regs_read_arr(270)(REG_OH_LINKS_OH10_VFAT8_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(8).sync_good;
    regs_read_arr(270)(REG_OH_LINKS_OH10_VFAT8_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT8_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(8).sync_error_cnt;
    regs_read_arr(270)(REG_OH_LINKS_OH10_VFAT8_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT8_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(8).daq_event_cnt;
    regs_read_arr(270)(REG_OH_LINKS_OH10_VFAT8_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT8_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(8).daq_crc_err_cnt;
    regs_read_arr(271)(REG_OH_LINKS_OH10_VFAT9_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(9).sync_good;
    regs_read_arr(271)(REG_OH_LINKS_OH10_VFAT9_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT9_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(9).sync_error_cnt;
    regs_read_arr(271)(REG_OH_LINKS_OH10_VFAT9_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT9_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(9).daq_event_cnt;
    regs_read_arr(271)(REG_OH_LINKS_OH10_VFAT9_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT9_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(9).daq_crc_err_cnt;
    regs_read_arr(272)(REG_OH_LINKS_OH10_VFAT10_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(10).sync_good;
    regs_read_arr(272)(REG_OH_LINKS_OH10_VFAT10_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT10_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(10).sync_error_cnt;
    regs_read_arr(272)(REG_OH_LINKS_OH10_VFAT10_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT10_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(10).daq_event_cnt;
    regs_read_arr(272)(REG_OH_LINKS_OH10_VFAT10_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT10_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(10).daq_crc_err_cnt;
    regs_read_arr(273)(REG_OH_LINKS_OH10_VFAT11_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(11).sync_good;
    regs_read_arr(273)(REG_OH_LINKS_OH10_VFAT11_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT11_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(11).sync_error_cnt;
    regs_read_arr(273)(REG_OH_LINKS_OH10_VFAT11_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT11_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(11).daq_event_cnt;
    regs_read_arr(273)(REG_OH_LINKS_OH10_VFAT11_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT11_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(11).daq_crc_err_cnt;
    regs_read_arr(274)(REG_OH_LINKS_OH10_VFAT12_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(12).sync_good;
    regs_read_arr(274)(REG_OH_LINKS_OH10_VFAT12_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT12_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(12).sync_error_cnt;
    regs_read_arr(274)(REG_OH_LINKS_OH10_VFAT12_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT12_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(12).daq_event_cnt;
    regs_read_arr(274)(REG_OH_LINKS_OH10_VFAT12_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT12_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(12).daq_crc_err_cnt;
    regs_read_arr(275)(REG_OH_LINKS_OH10_VFAT13_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(13).sync_good;
    regs_read_arr(275)(REG_OH_LINKS_OH10_VFAT13_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT13_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(13).sync_error_cnt;
    regs_read_arr(275)(REG_OH_LINKS_OH10_VFAT13_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT13_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(13).daq_event_cnt;
    regs_read_arr(275)(REG_OH_LINKS_OH10_VFAT13_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT13_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(13).daq_crc_err_cnt;
    regs_read_arr(276)(REG_OH_LINKS_OH10_VFAT14_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(14).sync_good;
    regs_read_arr(276)(REG_OH_LINKS_OH10_VFAT14_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT14_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(14).sync_error_cnt;
    regs_read_arr(276)(REG_OH_LINKS_OH10_VFAT14_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT14_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(14).daq_event_cnt;
    regs_read_arr(276)(REG_OH_LINKS_OH10_VFAT14_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT14_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(14).daq_crc_err_cnt;
    regs_read_arr(277)(REG_OH_LINKS_OH10_VFAT15_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(15).sync_good;
    regs_read_arr(277)(REG_OH_LINKS_OH10_VFAT15_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT15_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(15).sync_error_cnt;
    regs_read_arr(277)(REG_OH_LINKS_OH10_VFAT15_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT15_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(15).daq_event_cnt;
    regs_read_arr(277)(REG_OH_LINKS_OH10_VFAT15_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT15_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(15).daq_crc_err_cnt;
    regs_read_arr(278)(REG_OH_LINKS_OH10_VFAT16_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(16).sync_good;
    regs_read_arr(278)(REG_OH_LINKS_OH10_VFAT16_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT16_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(16).sync_error_cnt;
    regs_read_arr(278)(REG_OH_LINKS_OH10_VFAT16_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT16_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(16).daq_event_cnt;
    regs_read_arr(278)(REG_OH_LINKS_OH10_VFAT16_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT16_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(16).daq_crc_err_cnt;
    regs_read_arr(279)(REG_OH_LINKS_OH10_VFAT17_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(17).sync_good;
    regs_read_arr(279)(REG_OH_LINKS_OH10_VFAT17_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT17_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(17).sync_error_cnt;
    regs_read_arr(279)(REG_OH_LINKS_OH10_VFAT17_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT17_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(17).daq_event_cnt;
    regs_read_arr(279)(REG_OH_LINKS_OH10_VFAT17_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT17_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(17).daq_crc_err_cnt;
    regs_read_arr(280)(REG_OH_LINKS_OH10_VFAT18_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(18).sync_good;
    regs_read_arr(280)(REG_OH_LINKS_OH10_VFAT18_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT18_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(18).sync_error_cnt;
    regs_read_arr(280)(REG_OH_LINKS_OH10_VFAT18_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT18_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(18).daq_event_cnt;
    regs_read_arr(280)(REG_OH_LINKS_OH10_VFAT18_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT18_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(18).daq_crc_err_cnt;
    regs_read_arr(281)(REG_OH_LINKS_OH10_VFAT19_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(19).sync_good;
    regs_read_arr(281)(REG_OH_LINKS_OH10_VFAT19_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT19_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(19).sync_error_cnt;
    regs_read_arr(281)(REG_OH_LINKS_OH10_VFAT19_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT19_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(19).daq_event_cnt;
    regs_read_arr(281)(REG_OH_LINKS_OH10_VFAT19_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT19_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(19).daq_crc_err_cnt;
    regs_read_arr(282)(REG_OH_LINKS_OH10_VFAT20_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(20).sync_good;
    regs_read_arr(282)(REG_OH_LINKS_OH10_VFAT20_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT20_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(20).sync_error_cnt;
    regs_read_arr(282)(REG_OH_LINKS_OH10_VFAT20_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT20_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(20).daq_event_cnt;
    regs_read_arr(282)(REG_OH_LINKS_OH10_VFAT20_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT20_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(20).daq_crc_err_cnt;
    regs_read_arr(283)(REG_OH_LINKS_OH10_VFAT21_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(21).sync_good;
    regs_read_arr(283)(REG_OH_LINKS_OH10_VFAT21_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT21_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(21).sync_error_cnt;
    regs_read_arr(283)(REG_OH_LINKS_OH10_VFAT21_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT21_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(21).daq_event_cnt;
    regs_read_arr(283)(REG_OH_LINKS_OH10_VFAT21_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT21_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(21).daq_crc_err_cnt;
    regs_read_arr(284)(REG_OH_LINKS_OH10_VFAT22_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(22).sync_good;
    regs_read_arr(284)(REG_OH_LINKS_OH10_VFAT22_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT22_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(22).sync_error_cnt;
    regs_read_arr(284)(REG_OH_LINKS_OH10_VFAT22_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT22_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(22).daq_event_cnt;
    regs_read_arr(284)(REG_OH_LINKS_OH10_VFAT22_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT22_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(22).daq_crc_err_cnt;
    regs_read_arr(285)(REG_OH_LINKS_OH10_VFAT23_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(10)(23).sync_good;
    regs_read_arr(285)(REG_OH_LINKS_OH10_VFAT23_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT23_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(10)(23).sync_error_cnt;
    regs_read_arr(285)(REG_OH_LINKS_OH10_VFAT23_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH10_VFAT23_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(10)(23).daq_event_cnt;
    regs_read_arr(285)(REG_OH_LINKS_OH10_VFAT23_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH10_VFAT23_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(10)(23).daq_crc_err_cnt;
    regs_read_arr(286)(REG_OH_LINKS_OH11_GBT0_READY_BIT) <= gbt_link_status_arr_i(11 * g_NUM_GBTS_PER_OH + 0).gbt_rx_ready;
    regs_read_arr(286)(REG_OH_LINKS_OH11_GBT1_READY_BIT) <= gbt_link_status_arr_i(11 * g_NUM_GBTS_PER_OH + 1).gbt_rx_ready;
    regs_read_arr(286)(REG_OH_LINKS_OH11_GBT2_READY_BIT) <= gbt_link_status_arr_i(11 * g_NUM_GBTS_PER_OH + 2).gbt_rx_ready;
    regs_read_arr(286)(REG_OH_LINKS_OH11_GBT0_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(11 * g_NUM_GBTS_PER_OH + 0).gbt_rx_had_not_ready;
    regs_read_arr(286)(REG_OH_LINKS_OH11_GBT1_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(11 * g_NUM_GBTS_PER_OH + 1).gbt_rx_had_not_ready;
    regs_read_arr(286)(REG_OH_LINKS_OH11_GBT2_WAS_NOT_READY_BIT) <= gbt_link_status_arr_i(11 * g_NUM_GBTS_PER_OH + 2).gbt_rx_had_not_ready;
    regs_read_arr(286)(REG_OH_LINKS_OH11_GBT0_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(11 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_ovf;
    regs_read_arr(286)(REG_OH_LINKS_OH11_GBT1_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(11 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_ovf;
    regs_read_arr(286)(REG_OH_LINKS_OH11_GBT2_RX_HAD_OVERFLOW_BIT) <= gbt_link_status_arr_i(11 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_ovf;
    regs_read_arr(286)(REG_OH_LINKS_OH11_GBT0_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(11 * g_NUM_GBTS_PER_OH + 0).gbt_rx_sync_status.had_unf;
    regs_read_arr(286)(REG_OH_LINKS_OH11_GBT1_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(11 * g_NUM_GBTS_PER_OH + 1).gbt_rx_sync_status.had_unf;
    regs_read_arr(286)(REG_OH_LINKS_OH11_GBT2_RX_HAD_UNDERFLOW_BIT) <= gbt_link_status_arr_i(11 * g_NUM_GBTS_PER_OH + 2).gbt_rx_sync_status.had_unf;
    regs_read_arr(287)(REG_OH_LINKS_OH11_VFAT_MASK_MSB downto REG_OH_LINKS_OH11_VFAT_MASK_LSB) <= vfat_mask_arr(11);
    regs_read_arr(288)(REG_OH_LINKS_OH11_VFAT0_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(0).sync_good;
    regs_read_arr(288)(REG_OH_LINKS_OH11_VFAT0_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT0_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(0).sync_error_cnt;
    regs_read_arr(288)(REG_OH_LINKS_OH11_VFAT0_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT0_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(0).daq_event_cnt;
    regs_read_arr(288)(REG_OH_LINKS_OH11_VFAT0_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT0_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(0).daq_crc_err_cnt;
    regs_read_arr(289)(REG_OH_LINKS_OH11_VFAT1_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(1).sync_good;
    regs_read_arr(289)(REG_OH_LINKS_OH11_VFAT1_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT1_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(1).sync_error_cnt;
    regs_read_arr(289)(REG_OH_LINKS_OH11_VFAT1_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT1_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(1).daq_event_cnt;
    regs_read_arr(289)(REG_OH_LINKS_OH11_VFAT1_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT1_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(1).daq_crc_err_cnt;
    regs_read_arr(290)(REG_OH_LINKS_OH11_VFAT2_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(2).sync_good;
    regs_read_arr(290)(REG_OH_LINKS_OH11_VFAT2_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT2_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(2).sync_error_cnt;
    regs_read_arr(290)(REG_OH_LINKS_OH11_VFAT2_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT2_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(2).daq_event_cnt;
    regs_read_arr(290)(REG_OH_LINKS_OH11_VFAT2_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT2_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(2).daq_crc_err_cnt;
    regs_read_arr(291)(REG_OH_LINKS_OH11_VFAT3_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(3).sync_good;
    regs_read_arr(291)(REG_OH_LINKS_OH11_VFAT3_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT3_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(3).sync_error_cnt;
    regs_read_arr(291)(REG_OH_LINKS_OH11_VFAT3_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT3_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(3).daq_event_cnt;
    regs_read_arr(291)(REG_OH_LINKS_OH11_VFAT3_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT3_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(3).daq_crc_err_cnt;
    regs_read_arr(292)(REG_OH_LINKS_OH11_VFAT4_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(4).sync_good;
    regs_read_arr(292)(REG_OH_LINKS_OH11_VFAT4_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT4_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(4).sync_error_cnt;
    regs_read_arr(292)(REG_OH_LINKS_OH11_VFAT4_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT4_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(4).daq_event_cnt;
    regs_read_arr(292)(REG_OH_LINKS_OH11_VFAT4_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT4_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(4).daq_crc_err_cnt;
    regs_read_arr(293)(REG_OH_LINKS_OH11_VFAT5_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(5).sync_good;
    regs_read_arr(293)(REG_OH_LINKS_OH11_VFAT5_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT5_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(5).sync_error_cnt;
    regs_read_arr(293)(REG_OH_LINKS_OH11_VFAT5_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT5_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(5).daq_event_cnt;
    regs_read_arr(293)(REG_OH_LINKS_OH11_VFAT5_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT5_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(5).daq_crc_err_cnt;
    regs_read_arr(294)(REG_OH_LINKS_OH11_VFAT6_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(6).sync_good;
    regs_read_arr(294)(REG_OH_LINKS_OH11_VFAT6_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT6_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(6).sync_error_cnt;
    regs_read_arr(294)(REG_OH_LINKS_OH11_VFAT6_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT6_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(6).daq_event_cnt;
    regs_read_arr(294)(REG_OH_LINKS_OH11_VFAT6_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT6_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(6).daq_crc_err_cnt;
    regs_read_arr(295)(REG_OH_LINKS_OH11_VFAT7_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(7).sync_good;
    regs_read_arr(295)(REG_OH_LINKS_OH11_VFAT7_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT7_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(7).sync_error_cnt;
    regs_read_arr(295)(REG_OH_LINKS_OH11_VFAT7_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT7_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(7).daq_event_cnt;
    regs_read_arr(295)(REG_OH_LINKS_OH11_VFAT7_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT7_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(7).daq_crc_err_cnt;
    regs_read_arr(296)(REG_OH_LINKS_OH11_VFAT8_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(8).sync_good;
    regs_read_arr(296)(REG_OH_LINKS_OH11_VFAT8_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT8_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(8).sync_error_cnt;
    regs_read_arr(296)(REG_OH_LINKS_OH11_VFAT8_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT8_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(8).daq_event_cnt;
    regs_read_arr(296)(REG_OH_LINKS_OH11_VFAT8_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT8_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(8).daq_crc_err_cnt;
    regs_read_arr(297)(REG_OH_LINKS_OH11_VFAT9_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(9).sync_good;
    regs_read_arr(297)(REG_OH_LINKS_OH11_VFAT9_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT9_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(9).sync_error_cnt;
    regs_read_arr(297)(REG_OH_LINKS_OH11_VFAT9_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT9_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(9).daq_event_cnt;
    regs_read_arr(297)(REG_OH_LINKS_OH11_VFAT9_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT9_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(9).daq_crc_err_cnt;
    regs_read_arr(298)(REG_OH_LINKS_OH11_VFAT10_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(10).sync_good;
    regs_read_arr(298)(REG_OH_LINKS_OH11_VFAT10_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT10_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(10).sync_error_cnt;
    regs_read_arr(298)(REG_OH_LINKS_OH11_VFAT10_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT10_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(10).daq_event_cnt;
    regs_read_arr(298)(REG_OH_LINKS_OH11_VFAT10_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT10_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(10).daq_crc_err_cnt;
    regs_read_arr(299)(REG_OH_LINKS_OH11_VFAT11_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(11).sync_good;
    regs_read_arr(299)(REG_OH_LINKS_OH11_VFAT11_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT11_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(11).sync_error_cnt;
    regs_read_arr(299)(REG_OH_LINKS_OH11_VFAT11_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT11_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(11).daq_event_cnt;
    regs_read_arr(299)(REG_OH_LINKS_OH11_VFAT11_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT11_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(11).daq_crc_err_cnt;
    regs_read_arr(300)(REG_OH_LINKS_OH11_VFAT12_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(12).sync_good;
    regs_read_arr(300)(REG_OH_LINKS_OH11_VFAT12_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT12_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(12).sync_error_cnt;
    regs_read_arr(300)(REG_OH_LINKS_OH11_VFAT12_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT12_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(12).daq_event_cnt;
    regs_read_arr(300)(REG_OH_LINKS_OH11_VFAT12_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT12_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(12).daq_crc_err_cnt;
    regs_read_arr(301)(REG_OH_LINKS_OH11_VFAT13_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(13).sync_good;
    regs_read_arr(301)(REG_OH_LINKS_OH11_VFAT13_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT13_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(13).sync_error_cnt;
    regs_read_arr(301)(REG_OH_LINKS_OH11_VFAT13_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT13_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(13).daq_event_cnt;
    regs_read_arr(301)(REG_OH_LINKS_OH11_VFAT13_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT13_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(13).daq_crc_err_cnt;
    regs_read_arr(302)(REG_OH_LINKS_OH11_VFAT14_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(14).sync_good;
    regs_read_arr(302)(REG_OH_LINKS_OH11_VFAT14_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT14_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(14).sync_error_cnt;
    regs_read_arr(302)(REG_OH_LINKS_OH11_VFAT14_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT14_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(14).daq_event_cnt;
    regs_read_arr(302)(REG_OH_LINKS_OH11_VFAT14_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT14_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(14).daq_crc_err_cnt;
    regs_read_arr(303)(REG_OH_LINKS_OH11_VFAT15_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(15).sync_good;
    regs_read_arr(303)(REG_OH_LINKS_OH11_VFAT15_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT15_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(15).sync_error_cnt;
    regs_read_arr(303)(REG_OH_LINKS_OH11_VFAT15_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT15_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(15).daq_event_cnt;
    regs_read_arr(303)(REG_OH_LINKS_OH11_VFAT15_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT15_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(15).daq_crc_err_cnt;
    regs_read_arr(304)(REG_OH_LINKS_OH11_VFAT16_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(16).sync_good;
    regs_read_arr(304)(REG_OH_LINKS_OH11_VFAT16_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT16_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(16).sync_error_cnt;
    regs_read_arr(304)(REG_OH_LINKS_OH11_VFAT16_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT16_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(16).daq_event_cnt;
    regs_read_arr(304)(REG_OH_LINKS_OH11_VFAT16_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT16_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(16).daq_crc_err_cnt;
    regs_read_arr(305)(REG_OH_LINKS_OH11_VFAT17_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(17).sync_good;
    regs_read_arr(305)(REG_OH_LINKS_OH11_VFAT17_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT17_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(17).sync_error_cnt;
    regs_read_arr(305)(REG_OH_LINKS_OH11_VFAT17_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT17_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(17).daq_event_cnt;
    regs_read_arr(305)(REG_OH_LINKS_OH11_VFAT17_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT17_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(17).daq_crc_err_cnt;
    regs_read_arr(306)(REG_OH_LINKS_OH11_VFAT18_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(18).sync_good;
    regs_read_arr(306)(REG_OH_LINKS_OH11_VFAT18_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT18_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(18).sync_error_cnt;
    regs_read_arr(306)(REG_OH_LINKS_OH11_VFAT18_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT18_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(18).daq_event_cnt;
    regs_read_arr(306)(REG_OH_LINKS_OH11_VFAT18_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT18_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(18).daq_crc_err_cnt;
    regs_read_arr(307)(REG_OH_LINKS_OH11_VFAT19_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(19).sync_good;
    regs_read_arr(307)(REG_OH_LINKS_OH11_VFAT19_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT19_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(19).sync_error_cnt;
    regs_read_arr(307)(REG_OH_LINKS_OH11_VFAT19_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT19_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(19).daq_event_cnt;
    regs_read_arr(307)(REG_OH_LINKS_OH11_VFAT19_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT19_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(19).daq_crc_err_cnt;
    regs_read_arr(308)(REG_OH_LINKS_OH11_VFAT20_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(20).sync_good;
    regs_read_arr(308)(REG_OH_LINKS_OH11_VFAT20_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT20_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(20).sync_error_cnt;
    regs_read_arr(308)(REG_OH_LINKS_OH11_VFAT20_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT20_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(20).daq_event_cnt;
    regs_read_arr(308)(REG_OH_LINKS_OH11_VFAT20_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT20_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(20).daq_crc_err_cnt;
    regs_read_arr(309)(REG_OH_LINKS_OH11_VFAT21_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(21).sync_good;
    regs_read_arr(309)(REG_OH_LINKS_OH11_VFAT21_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT21_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(21).sync_error_cnt;
    regs_read_arr(309)(REG_OH_LINKS_OH11_VFAT21_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT21_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(21).daq_event_cnt;
    regs_read_arr(309)(REG_OH_LINKS_OH11_VFAT21_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT21_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(21).daq_crc_err_cnt;
    regs_read_arr(310)(REG_OH_LINKS_OH11_VFAT22_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(22).sync_good;
    regs_read_arr(310)(REG_OH_LINKS_OH11_VFAT22_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT22_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(22).sync_error_cnt;
    regs_read_arr(310)(REG_OH_LINKS_OH11_VFAT22_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT22_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(22).daq_event_cnt;
    regs_read_arr(310)(REG_OH_LINKS_OH11_VFAT22_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT22_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(22).daq_crc_err_cnt;
    regs_read_arr(311)(REG_OH_LINKS_OH11_VFAT23_LINK_GOOD_BIT) <= vfat3_link_status_arr_i(11)(23).sync_good;
    regs_read_arr(311)(REG_OH_LINKS_OH11_VFAT23_SYNC_ERR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT23_SYNC_ERR_CNT_LSB) <= vfat3_link_status_arr_i(11)(23).sync_error_cnt;
    regs_read_arr(311)(REG_OH_LINKS_OH11_VFAT23_DAQ_EVENT_CNT_MSB downto REG_OH_LINKS_OH11_VFAT23_DAQ_EVENT_CNT_LSB) <= vfat3_link_status_arr_i(11)(23).daq_event_cnt;
    regs_read_arr(311)(REG_OH_LINKS_OH11_VFAT23_DAQ_CRC_ERROR_CNT_MSB downto REG_OH_LINKS_OH11_VFAT23_DAQ_CRC_ERROR_CNT_LSB) <= vfat3_link_status_arr_i(11)(23).daq_crc_err_cnt;

    -- Connect write signals
    vfat_mask_arr(0) <= regs_write_arr(1)(REG_OH_LINKS_OH0_VFAT_MASK_MSB downto REG_OH_LINKS_OH0_VFAT_MASK_LSB);
    vfat_mask_arr(1) <= regs_write_arr(27)(REG_OH_LINKS_OH1_VFAT_MASK_MSB downto REG_OH_LINKS_OH1_VFAT_MASK_LSB);
    vfat_mask_arr(2) <= regs_write_arr(53)(REG_OH_LINKS_OH2_VFAT_MASK_MSB downto REG_OH_LINKS_OH2_VFAT_MASK_LSB);
    vfat_mask_arr(3) <= regs_write_arr(79)(REG_OH_LINKS_OH3_VFAT_MASK_MSB downto REG_OH_LINKS_OH3_VFAT_MASK_LSB);
    vfat_mask_arr(4) <= regs_write_arr(105)(REG_OH_LINKS_OH4_VFAT_MASK_MSB downto REG_OH_LINKS_OH4_VFAT_MASK_LSB);
    vfat_mask_arr(5) <= regs_write_arr(131)(REG_OH_LINKS_OH5_VFAT_MASK_MSB downto REG_OH_LINKS_OH5_VFAT_MASK_LSB);
    vfat_mask_arr(6) <= regs_write_arr(157)(REG_OH_LINKS_OH6_VFAT_MASK_MSB downto REG_OH_LINKS_OH6_VFAT_MASK_LSB);
    vfat_mask_arr(7) <= regs_write_arr(183)(REG_OH_LINKS_OH7_VFAT_MASK_MSB downto REG_OH_LINKS_OH7_VFAT_MASK_LSB);
    vfat_mask_arr(8) <= regs_write_arr(209)(REG_OH_LINKS_OH8_VFAT_MASK_MSB downto REG_OH_LINKS_OH8_VFAT_MASK_LSB);
    vfat_mask_arr(9) <= regs_write_arr(235)(REG_OH_LINKS_OH9_VFAT_MASK_MSB downto REG_OH_LINKS_OH9_VFAT_MASK_LSB);
    vfat_mask_arr(10) <= regs_write_arr(261)(REG_OH_LINKS_OH10_VFAT_MASK_MSB downto REG_OH_LINKS_OH10_VFAT_MASK_LSB);
    vfat_mask_arr(11) <= regs_write_arr(287)(REG_OH_LINKS_OH11_VFAT_MASK_MSB downto REG_OH_LINKS_OH11_VFAT_MASK_LSB);

    -- Connect write pulse signals

    -- Connect write done signals

    -- Connect read pulse signals

    -- Connect read ready signals

    -- Defaults
    regs_defaults(1)(REG_OH_LINKS_OH0_VFAT_MASK_MSB downto REG_OH_LINKS_OH0_VFAT_MASK_LSB) <= REG_OH_LINKS_OH0_VFAT_MASK_DEFAULT;
    regs_defaults(27)(REG_OH_LINKS_OH1_VFAT_MASK_MSB downto REG_OH_LINKS_OH1_VFAT_MASK_LSB) <= REG_OH_LINKS_OH1_VFAT_MASK_DEFAULT;
    regs_defaults(53)(REG_OH_LINKS_OH2_VFAT_MASK_MSB downto REG_OH_LINKS_OH2_VFAT_MASK_LSB) <= REG_OH_LINKS_OH2_VFAT_MASK_DEFAULT;
    regs_defaults(79)(REG_OH_LINKS_OH3_VFAT_MASK_MSB downto REG_OH_LINKS_OH3_VFAT_MASK_LSB) <= REG_OH_LINKS_OH3_VFAT_MASK_DEFAULT;
    regs_defaults(105)(REG_OH_LINKS_OH4_VFAT_MASK_MSB downto REG_OH_LINKS_OH4_VFAT_MASK_LSB) <= REG_OH_LINKS_OH4_VFAT_MASK_DEFAULT;
    regs_defaults(131)(REG_OH_LINKS_OH5_VFAT_MASK_MSB downto REG_OH_LINKS_OH5_VFAT_MASK_LSB) <= REG_OH_LINKS_OH5_VFAT_MASK_DEFAULT;
    regs_defaults(157)(REG_OH_LINKS_OH6_VFAT_MASK_MSB downto REG_OH_LINKS_OH6_VFAT_MASK_LSB) <= REG_OH_LINKS_OH6_VFAT_MASK_DEFAULT;
    regs_defaults(183)(REG_OH_LINKS_OH7_VFAT_MASK_MSB downto REG_OH_LINKS_OH7_VFAT_MASK_LSB) <= REG_OH_LINKS_OH7_VFAT_MASK_DEFAULT;
    regs_defaults(209)(REG_OH_LINKS_OH8_VFAT_MASK_MSB downto REG_OH_LINKS_OH8_VFAT_MASK_LSB) <= REG_OH_LINKS_OH8_VFAT_MASK_DEFAULT;
    regs_defaults(235)(REG_OH_LINKS_OH9_VFAT_MASK_MSB downto REG_OH_LINKS_OH9_VFAT_MASK_LSB) <= REG_OH_LINKS_OH9_VFAT_MASK_DEFAULT;
    regs_defaults(261)(REG_OH_LINKS_OH10_VFAT_MASK_MSB downto REG_OH_LINKS_OH10_VFAT_MASK_LSB) <= REG_OH_LINKS_OH10_VFAT_MASK_DEFAULT;
    regs_defaults(287)(REG_OH_LINKS_OH11_VFAT_MASK_MSB downto REG_OH_LINKS_OH11_VFAT_MASK_LSB) <= REG_OH_LINKS_OH11_VFAT_MASK_DEFAULT;

    -- Define writable regs
    regs_writable_arr(1) <= '1';
    regs_writable_arr(27) <= '1';
    regs_writable_arr(53) <= '1';
    regs_writable_arr(79) <= '1';
    regs_writable_arr(105) <= '1';
    regs_writable_arr(131) <= '1';
    regs_writable_arr(157) <= '1';
    regs_writable_arr(183) <= '1';
    regs_writable_arr(209) <= '1';
    regs_writable_arr(235) <= '1';
    regs_writable_arr(261) <= '1';
    regs_writable_arr(287) <= '1';

    --==== Registers end ============================================================================
    
end oh_link_regs_arch;

